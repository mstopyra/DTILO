magic
tech sky130A
timestamp 1702609360
<< nmos >>
rect 2600 14500 3000 17700
rect 12100 14500 12500 17700
rect 13600 14500 14000 17700
rect 2600 10900 3000 14100
rect 12300 10800 12700 14000
<< ndiff >>
rect 2300 17500 2600 17700
rect 2300 14700 2400 17500
rect 2500 14700 2600 17500
rect 2300 14500 2600 14700
rect 3000 17500 3300 17700
rect 3000 14700 3100 17500
rect 3200 14700 3300 17500
rect 3000 14500 3300 14700
rect 11800 17500 12100 17700
rect 11800 14700 11900 17500
rect 12000 14700 12100 17500
rect 11800 14500 12100 14700
rect 12500 17500 12800 17700
rect 12500 14700 12600 17500
rect 12700 14700 12800 17500
rect 12500 14500 12800 14700
rect 13300 17500 13600 17700
rect 13300 14700 13400 17500
rect 13500 14700 13600 17500
rect 13300 14500 13600 14700
rect 14000 17500 14300 17700
rect 14000 14700 14100 17500
rect 14200 14700 14300 17500
rect 14000 14500 14300 14700
rect 2300 13900 2600 14100
rect 2300 11100 2400 13900
rect 2500 11100 2600 13900
rect 2300 10900 2600 11100
rect 3000 13900 3300 14100
rect 3000 11100 3100 13900
rect 3200 11100 3300 13900
rect 3000 10900 3300 11100
rect 12000 13800 12300 14000
rect 12000 11000 12100 13800
rect 12200 11000 12300 13800
rect 12000 10800 12300 11000
rect 12700 13800 13000 14000
rect 12700 11000 12800 13800
rect 12900 11000 13000 13800
rect 12700 10800 13000 11000
<< ndiffc >>
rect 2400 14700 2500 17500
rect 3100 14700 3200 17500
rect 11900 14700 12000 17500
rect 12600 14700 12700 17500
rect 13400 14700 13500 17500
rect 14100 14700 14200 17500
rect 2400 11100 2500 13900
rect 3100 11100 3200 13900
rect 12100 11000 12200 13800
rect 12800 11000 12900 13800
<< psubdiff >>
rect 2000 17500 2300 17700
rect 2000 16210 2100 17500
rect 2002 15948 2100 16210
rect 2000 14700 2100 15948
rect 2200 14700 2300 17500
rect 2000 14500 2300 14700
rect 11530 17600 11800 17700
rect 11530 14600 11600 17600
rect 11700 14600 11800 17600
rect 11530 14500 11800 14600
rect 13000 17500 13300 17700
rect 13000 14700 13100 17500
rect 13200 14700 13300 17500
rect 13000 14500 13300 14700
rect 2000 13900 2300 14100
rect 2000 11100 2100 13900
rect 2200 11100 2300 13900
rect 2000 10900 2300 11100
rect 11700 13800 12000 14000
rect 11700 11000 11800 13800
rect 11900 11000 12000 13800
rect 11700 10800 12000 11000
<< psubdiffcont >>
rect 2100 14700 2200 17500
rect 11600 14600 11700 17600
rect 13100 14700 13200 17500
rect 2100 11100 2200 13900
rect 11800 11000 11900 13800
<< poly >>
rect 11200 17950 12500 18000
rect 11200 17850 12150 17950
rect 12450 17850 12500 17950
rect 11200 17800 12500 17850
rect 13200 17950 14000 18000
rect 13200 17850 13250 17950
rect 13450 17850 14000 17950
rect 13200 17800 14000 17850
rect 2600 17700 3000 17800
rect 12100 17700 12500 17800
rect 13600 17700 14000 17800
rect 2600 14350 3000 14500
rect 12100 14400 12500 14500
rect 2600 14250 2650 14350
rect 2950 14250 3000 14350
rect 13600 14300 14000 14500
rect 2600 14100 3000 14250
rect 12300 14100 14000 14300
rect 12300 14000 12700 14100
rect 2600 10800 3000 10900
rect 12300 10700 12700 10800
<< polycont >>
rect 12150 17850 12450 17950
rect 13250 17850 13450 17950
rect 2650 14250 2950 14350
<< locali >>
rect 11600 17600 11700 18000
rect 12100 17950 12500 18000
rect 12100 17850 12150 17950
rect 12450 17850 12500 17950
rect 12100 17800 12500 17850
rect 13200 17950 13500 18000
rect 13200 17850 13250 17950
rect 13450 17850 13500 17950
rect 13200 17600 13500 17850
rect 2000 17500 2600 17600
rect 2000 16210 2100 17500
rect 2002 15948 2100 16210
rect 2000 14700 2100 15948
rect 2200 14700 2400 17500
rect 2500 14700 2600 17500
rect 2000 14600 2600 14700
rect 3000 17500 3300 17600
rect 3000 14700 3100 17500
rect 3200 14700 3300 17500
rect 3000 14600 3300 14700
rect 11800 17500 12100 17600
rect 11800 14700 11900 17500
rect 12000 14700 12100 17500
rect 11800 14600 12100 14700
rect 12500 17500 12800 17600
rect 12500 14700 12600 17500
rect 12700 14700 12800 17500
rect 12500 14600 12800 14700
rect 13000 17500 13600 17600
rect 13000 14700 13100 17500
rect 13200 14700 13400 17500
rect 13500 14700 13600 17500
rect 13000 14600 13600 14700
rect 14000 17500 14300 17600
rect 14000 14700 14100 17500
rect 14200 14700 14300 17500
rect 14000 14600 14300 14700
rect 2400 14400 2500 14600
rect 2400 14350 3000 14400
rect 2400 14250 2650 14350
rect 2950 14250 3000 14350
rect 2400 14200 3000 14250
rect 11600 14300 11700 14600
rect 12500 14500 12700 14600
rect 14000 14500 14200 14600
rect 11600 14200 11900 14300
rect 2400 14000 2500 14200
rect 2000 13900 2600 14000
rect 2000 11100 2100 13900
rect 2200 11100 2400 13900
rect 2500 11100 2600 13900
rect 2000 11000 2600 11100
rect 3000 13900 3300 14000
rect 11800 13900 11900 14200
rect 3000 11100 3100 13900
rect 3200 11100 3300 13900
rect 3000 11000 3300 11100
rect 11700 13800 12300 13900
rect 11700 11000 11800 13800
rect 11900 11000 12100 13800
rect 12200 11000 12300 13800
rect 11200 10900 11500 11000
rect 11700 10900 12300 11000
rect 12700 13800 13000 13900
rect 12700 11000 12800 13800
rect 12900 11000 13000 13800
rect 12700 10900 13000 11000
rect 11300 10700 11500 10900
rect 12700 10800 12900 10900
rect 11250 10650 11450 10700
rect 11250 10500 11300 10650
rect 11400 10600 11450 10650
<< viali >>
rect 2400 14700 2500 17500
rect 3100 16000 3200 16200
rect 11900 16000 12000 16200
rect 12600 15000 12700 15200
rect 13400 14700 13500 17500
rect 14100 15950 14200 16250
rect 2400 11100 2500 13900
rect 3100 12200 3200 12400
rect 12100 11000 12200 13800
rect 12800 12150 12900 12450
rect 11300 10550 11400 10650
<< metal1 >>
rect 2300 17500 2600 17600
rect 2300 14700 2400 17500
rect 2500 14700 2600 17500
rect 13300 17500 13600 17600
rect 13300 16300 13400 17500
rect 3050 16200 3500 16300
rect 3050 16000 3100 16200
rect 3200 16000 3500 16200
rect 3050 15900 3500 16000
rect 11500 16200 12400 16300
rect 11500 16000 11900 16200
rect 12000 16000 12400 16200
rect 11500 15900 12400 16000
rect 13000 15900 13400 16300
rect 12500 15200 12800 15300
rect 12500 15000 12600 15200
rect 12700 15000 12800 15200
rect 12500 14900 12800 15000
rect 2300 13900 2600 14700
rect 13300 14700 13400 15900
rect 13500 14700 13600 17500
rect 14000 16250 14250 16300
rect 14000 15950 14100 16250
rect 14200 15950 14250 16250
rect 14000 15900 14250 15950
rect 13300 14500 13600 14700
rect 2300 11100 2400 13900
rect 2500 11100 2600 13900
rect 12000 14100 13600 14500
rect 12000 13800 12700 14100
rect 3000 12400 3500 12500
rect 3000 12200 3100 12400
rect 3200 12200 3500 12400
rect 3000 12100 3500 12200
rect 11500 12450 11700 12500
rect 11500 12150 11550 12450
rect 11650 12150 11700 12450
rect 11500 12100 11700 12150
rect 2300 10000 2600 11100
rect 12000 11000 12100 13800
rect 12200 11000 12700 13800
rect 12750 12450 12950 12500
rect 12750 12150 12800 12450
rect 12900 12150 12950 12450
rect 12750 12100 12950 12150
rect 11250 10650 11300 10700
rect 11000 10550 11300 10650
rect 11250 10500 11300 10550
rect 12000 10000 12700 11000
rect 2300 6800 3500 10000
rect 11500 6800 12700 10000
<< via1 >>
rect 3100 16000 3200 16200
rect 11900 16000 12000 16200
rect 12600 15000 12700 15200
rect 14100 15950 14200 16250
rect 3100 12200 3200 12400
rect 11550 12150 11650 12450
rect 12800 12150 12900 12450
rect 11300 10550 11400 10650
<< metal2 >>
rect 2000 16210 3300 16300
rect 2002 16200 3300 16210
rect 2002 16000 3100 16200
rect 3200 16000 3300 16200
rect 2002 15948 3300 16000
rect 2000 15900 3300 15948
rect 11800 16250 14250 16300
rect 11800 16200 14100 16250
rect 11800 16000 11900 16200
rect 12000 16000 14100 16200
rect 11800 15950 14100 16000
rect 14200 15950 14250 16250
rect 11800 15900 14250 15950
rect 11100 15200 14900 15300
rect 11100 15000 12600 15200
rect 12700 15000 14900 15200
rect 11100 14900 14900 15000
rect 2000 12400 3300 12500
rect 2000 12200 3100 12400
rect 3200 12200 3300 12400
rect 2000 12100 3300 12200
rect 11100 10700 11400 14900
rect 11500 12450 14900 12500
rect 11500 12150 11550 12450
rect 11650 12150 12800 12450
rect 12900 12150 14900 12450
rect 11500 12100 14900 12150
rect 11250 10650 11450 10700
rect 11250 10550 11300 10650
rect 11400 10550 11450 10650
rect 11250 10500 11450 10550
use DAC_block  DAC_block_14
timestamp 1702609360
transform 1 0 1800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_15
timestamp 1702609360
transform 1 0 7800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_16
timestamp 1702609360
transform 1 0 3800 0 1 10700
box 1700 -10800 3700 7300
use DAC_block  DAC_block_20
timestamp 1702609360
transform 1 0 5800 0 1 10700
box 1700 -10800 3700 7300
<< labels >>
flabel metal2 2000 12300 2000 12300 0 FreeSans 800 0 0 0 I_OUT
port 3 nsew
flabel metal1 2300 8300 2300 8300 0 FreeSans 800 0 0 0 VN
port 16 nsew
flabel space 3500 3300 3500 3300 0 FreeSans 800 0 0 0 VP
port 18 nsew
flabel space 8800 -100 8800 -100 0 FreeSans 800 0 0 0 D_1
port 10 nsew
flabel space 10800 -100 10800 -100 0 FreeSans 800 0 0 0 D_0
port 11 nsew
flabel metal2 14900 12300 14900 12300 0 FreeSans 800 0 0 0 I_OUT_LD
port 14 nsew
flabel metal2 14900 15100 14900 15100 0 FreeSans 800 0 0 0 I_DUMP
port 12 nsew
flabel space 6800 -100 6800 -100 0 FreeSans 800 0 0 0 D_2
port 6 nsew
flabel space 4800 -100 4800 -100 0 FreeSans 800 0 0 0 D_3
port 5 nsew
flabel space 3500 17900 3500 17900 0 FreeSans 800 0 0 0 VDD
port 19 nsew
<< end >>

magic
tech sky130A
timestamp 1702606600
<< nwell >>
rect 695 965 1115 1500
<< nmos >>
rect 775 705 790 805
rect 860 705 875 805
rect 775 405 790 505
rect 860 405 875 505
rect 940 405 955 805
rect 1030 705 1045 805
rect 1030 405 1045 505
<< pmos >>
rect 765 1290 780 1390
rect 830 1290 845 1390
rect 765 1020 780 1120
rect 830 1020 845 1120
rect 935 990 950 1390
rect 1010 1290 1025 1390
rect 1010 990 1025 1090
<< ndiff >>
rect 725 790 775 805
rect 725 720 740 790
rect 760 720 775 790
rect 725 705 775 720
rect 790 790 860 805
rect 790 720 825 790
rect 845 720 860 790
rect 790 705 860 720
rect 875 705 940 805
rect 915 505 940 705
rect 725 490 775 505
rect 725 420 740 490
rect 760 420 775 490
rect 725 405 775 420
rect 790 490 860 505
rect 790 420 825 490
rect 845 420 860 490
rect 790 405 860 420
rect 875 405 940 505
rect 955 790 1030 805
rect 955 720 970 790
rect 990 720 1030 790
rect 955 705 1030 720
rect 1045 790 1095 805
rect 1045 720 1060 790
rect 1080 720 1095 790
rect 1045 705 1095 720
rect 955 505 980 705
rect 955 490 1030 505
rect 955 420 970 490
rect 990 420 1030 490
rect 955 405 1030 420
rect 1045 490 1096 505
rect 1045 420 1060 490
rect 1080 420 1096 490
rect 1045 405 1096 420
<< pdiff >>
rect 715 1375 765 1390
rect 715 1305 730 1375
rect 750 1305 765 1375
rect 715 1290 765 1305
rect 780 1375 830 1390
rect 780 1305 795 1375
rect 815 1305 830 1375
rect 780 1290 830 1305
rect 845 1375 935 1390
rect 845 1290 900 1375
rect 885 1120 900 1290
rect 715 1105 765 1120
rect 715 1035 730 1105
rect 750 1035 765 1105
rect 715 1020 765 1035
rect 780 1105 830 1120
rect 780 1035 795 1105
rect 815 1035 830 1105
rect 780 1020 830 1035
rect 845 1020 900 1120
rect 885 1005 900 1020
rect 920 1005 935 1375
rect 885 990 935 1005
rect 950 1290 1010 1390
rect 1025 1375 1080 1390
rect 1025 1305 1045 1375
rect 1065 1305 1080 1375
rect 1025 1290 1080 1305
rect 950 1090 1000 1290
rect 950 990 1010 1090
rect 1025 1075 1075 1090
rect 1025 1005 1040 1075
rect 1060 1005 1075 1075
rect 1025 990 1075 1005
<< ndiffc >>
rect 740 720 760 790
rect 825 720 845 790
rect 740 420 760 490
rect 825 420 845 490
rect 970 720 990 790
rect 1060 720 1080 790
rect 970 420 990 490
rect 1060 420 1080 490
<< pdiffc >>
rect 730 1305 750 1375
rect 795 1305 815 1375
rect 730 1035 750 1105
rect 795 1035 815 1105
rect 900 1005 920 1375
rect 1045 1305 1065 1375
rect 1040 1005 1060 1075
<< psubdiff >>
rect 775 340 975 355
rect 775 315 790 340
rect 960 315 975 340
rect 775 300 975 315
<< nsubdiff >>
rect 970 1460 1070 1475
rect 970 1440 985 1460
rect 1055 1440 1070 1460
rect 970 1425 1070 1440
<< psubdiffcont >>
rect 790 315 960 340
<< nsubdiffcont >>
rect 985 1440 1055 1460
<< poly >>
rect 735 1445 780 1450
rect 735 1440 950 1445
rect 735 1415 745 1440
rect 770 1430 950 1440
rect 770 1415 780 1430
rect 735 1405 780 1415
rect 765 1390 780 1405
rect 830 1390 845 1405
rect 935 1390 950 1430
rect 1010 1390 1025 1405
rect 765 1275 780 1290
rect 830 1245 845 1290
rect 785 1230 845 1245
rect 785 1220 800 1230
rect 755 1210 800 1220
rect 755 1185 765 1210
rect 790 1185 800 1210
rect 755 1175 800 1185
rect 825 1170 870 1180
rect 825 1145 835 1170
rect 860 1145 870 1170
rect 825 1135 870 1145
rect 765 1120 780 1135
rect 830 1120 845 1135
rect 765 945 780 1020
rect 830 980 845 1020
rect 1010 1190 1025 1290
rect 1050 1265 1095 1275
rect 1050 1240 1060 1265
rect 1085 1245 1095 1265
rect 1085 1240 1100 1245
rect 1050 1230 1100 1240
rect 1010 1180 1060 1190
rect 1010 1155 1025 1180
rect 1050 1155 1060 1180
rect 1010 1145 1060 1155
rect 1085 1120 1100 1230
rect 1010 1105 1100 1120
rect 1010 1090 1025 1105
rect 830 965 875 980
rect 735 935 780 945
rect 735 910 745 935
rect 770 910 780 935
rect 735 900 780 910
rect 775 805 790 820
rect 860 805 875 965
rect 935 940 950 990
rect 1010 955 1025 990
rect 1005 940 1025 955
rect 905 930 950 940
rect 905 905 915 930
rect 940 905 950 930
rect 905 895 950 905
rect 975 930 1020 940
rect 975 905 985 930
rect 1010 905 1020 930
rect 975 895 1020 905
rect 1050 930 1095 940
rect 1050 905 1060 930
rect 1085 905 1095 930
rect 1050 895 1095 905
rect 925 870 940 895
rect 925 855 955 870
rect 940 805 955 855
rect 1055 835 1070 895
rect 1030 820 1070 835
rect 1030 805 1045 820
rect 775 690 790 705
rect 860 690 875 705
rect 750 680 795 690
rect 750 655 760 680
rect 785 655 795 680
rect 750 645 795 655
rect 855 680 900 690
rect 855 655 865 680
rect 890 655 900 680
rect 855 645 900 655
rect 705 610 750 620
rect 705 585 715 610
rect 740 585 750 610
rect 705 575 750 585
rect 775 505 790 645
rect 830 600 875 610
rect 830 575 840 600
rect 865 575 875 600
rect 830 565 875 575
rect 860 505 875 565
rect 1030 695 1045 705
rect 1020 690 1045 695
rect 990 680 1045 690
rect 990 655 1000 680
rect 1025 655 1035 680
rect 990 645 1035 655
rect 1030 600 1075 610
rect 1030 575 1040 600
rect 1065 575 1075 600
rect 1030 565 1075 575
rect 1030 505 1045 565
rect 775 390 790 405
rect 860 390 875 405
rect 940 390 955 405
rect 1030 390 1045 405
rect 1000 380 1045 390
rect 1000 355 1010 380
rect 1035 355 1045 380
rect 1000 345 1045 355
<< polycont >>
rect 745 1415 770 1440
rect 765 1185 790 1210
rect 835 1145 860 1170
rect 1060 1240 1085 1265
rect 1025 1155 1050 1180
rect 745 910 770 935
rect 915 905 940 930
rect 985 905 1010 930
rect 1060 905 1085 930
rect 760 655 785 680
rect 865 655 890 680
rect 715 585 740 610
rect 840 575 865 600
rect 1000 655 1025 680
rect 1040 575 1065 600
rect 1010 355 1035 380
<< locali >>
rect 975 1460 1065 1470
rect 735 1440 780 1450
rect 735 1415 745 1440
rect 770 1415 780 1440
rect 975 1440 985 1460
rect 1055 1440 1065 1460
rect 975 1430 1065 1440
rect 735 1405 780 1415
rect 720 1375 760 1385
rect 720 1345 730 1375
rect 695 1325 730 1345
rect 720 1305 730 1325
rect 750 1305 760 1375
rect 720 1295 760 1305
rect 785 1375 825 1385
rect 785 1305 795 1375
rect 815 1305 825 1375
rect 785 1295 825 1305
rect 890 1375 930 1385
rect 800 1275 820 1295
rect 800 1255 870 1275
rect 755 1210 800 1220
rect 755 1185 765 1210
rect 790 1195 800 1210
rect 790 1185 805 1195
rect 755 1175 805 1185
rect 850 1180 870 1255
rect 785 1115 805 1175
rect 825 1170 870 1180
rect 825 1145 835 1170
rect 860 1145 870 1170
rect 825 1135 870 1145
rect 720 1105 760 1115
rect 720 1075 730 1105
rect 695 1055 730 1075
rect 720 1035 730 1055
rect 750 1035 760 1105
rect 720 1025 760 1035
rect 785 1105 825 1115
rect 785 1035 795 1105
rect 815 1050 825 1105
rect 815 1035 835 1050
rect 785 1025 835 1035
rect 735 935 780 945
rect 735 910 745 935
rect 770 910 780 935
rect 735 900 780 910
rect 815 800 835 1025
rect 890 1005 900 1375
rect 920 1005 930 1375
rect 1035 1375 1075 1385
rect 1035 1305 1045 1375
rect 1065 1345 1075 1375
rect 1065 1325 1115 1345
rect 1065 1305 1075 1325
rect 1035 1295 1075 1305
rect 1050 1275 1070 1295
rect 1050 1265 1095 1275
rect 1050 1240 1060 1265
rect 1085 1240 1095 1265
rect 1050 1230 1095 1240
rect 1015 1180 1060 1190
rect 1015 1155 1025 1180
rect 1050 1155 1060 1180
rect 1015 1145 1060 1155
rect 1015 1085 1035 1145
rect 1015 1075 1070 1085
rect 1015 1060 1040 1075
rect 890 995 930 1005
rect 1030 1005 1040 1060
rect 1060 1055 1115 1075
rect 1060 1005 1070 1055
rect 1030 995 1070 1005
rect 1050 940 1070 995
rect 905 930 950 940
rect 905 905 915 930
rect 940 905 950 930
rect 905 895 950 905
rect 975 930 1020 940
rect 975 905 985 930
rect 1010 905 1020 930
rect 975 895 1020 905
rect 1050 930 1095 940
rect 1050 905 1060 930
rect 1085 905 1095 930
rect 1050 895 1095 905
rect 990 840 1010 895
rect 990 820 1090 840
rect 1070 800 1090 820
rect 730 790 770 800
rect 730 750 740 790
rect 710 720 740 750
rect 760 720 770 790
rect 710 710 770 720
rect 815 790 855 800
rect 815 720 825 790
rect 845 720 855 790
rect 815 710 855 720
rect 960 790 1000 800
rect 960 720 970 790
rect 990 720 1000 790
rect 960 710 1000 720
rect 1050 790 1090 800
rect 1050 720 1060 790
rect 1080 720 1090 790
rect 1050 710 1090 720
rect 710 620 730 710
rect 750 680 795 690
rect 750 655 760 680
rect 785 655 795 680
rect 750 645 795 655
rect 705 610 750 620
rect 705 585 715 610
rect 740 585 750 610
rect 815 610 835 710
rect 855 680 900 690
rect 855 655 865 680
rect 890 665 900 680
rect 990 680 1035 690
rect 890 655 915 665
rect 855 645 915 655
rect 815 600 875 610
rect 815 585 840 600
rect 705 575 750 585
rect 830 575 840 585
rect 865 575 875 600
rect 830 565 875 575
rect 895 545 915 645
rect 835 525 915 545
rect 990 655 1000 680
rect 1025 655 1035 680
rect 990 645 1035 655
rect 990 545 1010 645
rect 1070 610 1090 710
rect 1030 600 1090 610
rect 1030 575 1040 600
rect 1065 590 1090 600
rect 1065 575 1075 590
rect 1030 565 1075 575
rect 990 525 1070 545
rect 835 500 855 525
rect 1050 500 1070 525
rect 730 490 770 500
rect 730 420 740 490
rect 760 420 770 490
rect 730 410 770 420
rect 815 490 855 500
rect 815 420 825 490
rect 845 420 855 490
rect 815 410 855 420
rect 960 490 1000 500
rect 960 420 970 490
rect 990 420 1000 490
rect 960 410 1000 420
rect 1050 490 1090 500
rect 1050 420 1060 490
rect 1080 420 1090 490
rect 1050 410 1090 420
rect 740 390 760 410
rect 740 380 1045 390
rect 740 370 1010 380
rect 1000 355 1010 370
rect 1035 355 1045 380
rect 780 340 970 350
rect 1000 345 1045 355
rect 780 315 790 340
rect 960 315 970 340
rect 780 305 970 315
<< viali >>
rect 745 1415 770 1440
rect 985 1440 1055 1460
rect 745 910 770 935
rect 900 1005 920 1375
rect 915 905 940 930
rect 760 655 785 680
rect 715 585 740 610
rect 1000 655 1025 680
rect 970 420 990 490
rect 790 315 960 340
<< metal1 >>
rect 695 1465 1115 1500
rect 845 1460 1105 1465
rect 735 1440 780 1450
rect 735 1415 745 1440
rect 770 1415 780 1440
rect 735 940 780 1415
rect 845 1440 985 1460
rect 1055 1440 1105 1460
rect 845 1375 1105 1440
rect 845 1005 900 1375
rect 920 1005 1105 1375
rect 845 985 1105 1005
rect 695 935 1115 940
rect 695 910 745 935
rect 770 930 1115 935
rect 770 910 915 930
rect 695 905 915 910
rect 940 905 1115 930
rect 695 895 1115 905
rect 765 690 780 895
rect 750 680 795 690
rect 750 655 760 680
rect 785 655 795 680
rect 990 680 1035 690
rect 990 675 1000 680
rect 750 645 795 655
rect 865 660 1000 675
rect 705 610 750 620
rect 705 585 715 610
rect 740 605 750 610
rect 865 605 880 660
rect 990 655 1000 660
rect 1025 655 1035 680
rect 990 645 1035 655
rect 740 590 880 605
rect 740 585 750 590
rect 705 575 750 585
rect 695 490 1115 505
rect 695 420 970 490
rect 990 420 1115 490
rect 695 405 1115 420
rect 770 340 980 405
rect 770 315 790 340
rect 960 315 980 340
rect 770 295 980 315
<< labels >>
rlabel locali 1115 1335 1115 1335 3 Q_NOT
rlabel locali 1115 1065 1115 1065 3 Q
rlabel locali 695 1065 695 1065 7 D
rlabel locali 695 1335 695 1335 7 D_NOT
rlabel metal1 695 1485 695 1485 7 IN_RO
port 1 w
rlabel metal1 695 430 695 430 7 GND
port 3 w
rlabel metal1 695 920 695 920 7 IN_RO
<< end >>

magic
tech sky130A
timestamp 1702260771
<< nwell >>
rect -650 -200 13550 3350
rect -650 -250 13500 -200
<< nmos >>
rect -100 -3800 300 -600
rect 1050 -3800 1450 -600
rect 1700 -3800 2100 -600
rect 3100 -3800 3500 -600
rect 3750 -3800 4150 -600
rect 5150 -3800 5550 -600
rect 5600 -3800 6000 -600
rect 6900 -3800 7300 -600
rect 7350 -3800 7750 -600
rect 8750 -3800 9150 -600
rect 9400 -3800 9800 -600
rect 10800 -3800 11200 -600
rect 11450 -3800 11850 -600
rect 12600 -3800 13000 -600
<< pmos >>
rect -100 -50 300 3150
rect 1050 -50 1450 3150
rect 1500 -50 1900 3150
rect 3150 -50 3550 3150
rect 3600 -50 4000 3150
rect 5150 -50 5550 3150
rect 5600 -50 6000 3150
rect 6900 -50 7300 3150
rect 7350 -50 7750 3150
rect 8900 -50 9300 3150
rect 9350 -50 9750 3150
rect 11000 -50 11400 3150
rect 11450 -50 11850 3150
rect 12600 -50 13000 3150
<< ndiff >>
rect -350 -700 -100 -600
rect -350 -3700 -250 -700
rect -200 -3700 -100 -700
rect -350 -3800 -100 -3700
rect 300 -700 550 -600
rect 800 -700 1050 -600
rect 300 -3700 400 -700
rect 450 -3700 550 -700
rect 800 -3700 900 -700
rect 950 -3700 1050 -700
rect 300 -3800 550 -3700
rect 800 -3800 1050 -3700
rect 1450 -700 1700 -600
rect 1450 -3700 1550 -700
rect 1600 -3700 1700 -700
rect 1450 -3800 1700 -3700
rect 2100 -700 2350 -600
rect 2100 -3700 2200 -700
rect 2250 -3700 2350 -700
rect 2100 -3800 2350 -3700
rect 2850 -700 3100 -600
rect 2850 -3700 2950 -700
rect 3000 -3700 3100 -700
rect 2850 -3800 3100 -3700
rect 3500 -700 3750 -600
rect 3500 -3700 3600 -700
rect 3650 -3700 3750 -700
rect 3500 -3800 3750 -3700
rect 4150 -700 4400 -600
rect 4150 -3700 4250 -700
rect 4300 -3700 4400 -700
rect 4150 -3800 4400 -3700
rect 4900 -700 5150 -600
rect 4900 -3700 5000 -700
rect 5050 -3700 5150 -700
rect 4900 -3800 5150 -3700
rect 5550 -3800 5600 -600
rect 6000 -700 6250 -600
rect 6000 -3700 6100 -700
rect 6150 -3700 6250 -700
rect 6000 -3800 6250 -3700
rect 6650 -700 6900 -600
rect 6650 -3700 6750 -700
rect 6800 -3700 6900 -700
rect 6650 -3800 6900 -3700
rect 7300 -3800 7350 -600
rect 7750 -700 8000 -600
rect 7750 -3700 7850 -700
rect 7900 -3700 8000 -700
rect 7750 -3800 8000 -3700
rect 8500 -700 8750 -600
rect 8500 -3700 8600 -700
rect 8650 -3700 8750 -700
rect 8500 -3800 8750 -3700
rect 9150 -700 9400 -600
rect 9150 -3700 9250 -700
rect 9300 -3700 9400 -700
rect 9150 -3800 9400 -3700
rect 9800 -700 10050 -600
rect 9800 -3700 9900 -700
rect 9950 -3700 10050 -700
rect 9800 -3800 10050 -3700
rect 10550 -700 10800 -600
rect 10550 -3700 10650 -700
rect 10700 -3700 10800 -700
rect 10550 -3800 10800 -3700
rect 11200 -700 11450 -600
rect 11200 -3700 11300 -700
rect 11350 -3700 11450 -700
rect 11200 -3800 11450 -3700
rect 11850 -700 12100 -600
rect 12350 -700 12600 -600
rect 11850 -3700 11950 -700
rect 12000 -3700 12100 -700
rect 12350 -3700 12450 -700
rect 12500 -3700 12600 -700
rect 11850 -3800 12100 -3700
rect 12350 -3800 12600 -3700
rect 13000 -700 13250 -600
rect 13000 -3700 13100 -700
rect 13150 -3700 13250 -700
rect 13000 -3800 13250 -3700
<< pdiff >>
rect -350 3050 -100 3150
rect -350 50 -250 3050
rect -200 50 -100 3050
rect -350 -50 -100 50
rect 300 3050 550 3150
rect 800 3050 1050 3150
rect 300 50 400 3050
rect 450 50 550 3050
rect 800 50 900 3050
rect 950 50 1050 3050
rect 300 -50 550 50
rect 800 -50 1050 50
rect 1450 -50 1500 3150
rect 1900 3050 2150 3150
rect 1900 50 2000 3050
rect 2050 50 2150 3050
rect 1900 -50 2150 50
rect 2900 3050 3150 3150
rect 2900 50 3000 3050
rect 3050 50 3150 3050
rect 2900 -50 3150 50
rect 3550 -50 3600 3150
rect 4000 3050 4250 3150
rect 4000 50 4100 3050
rect 4150 50 4250 3050
rect 4000 -50 4250 50
rect 4900 3050 5150 3150
rect 4900 50 5000 3050
rect 5050 50 5150 3050
rect 4900 -50 5150 50
rect 5550 -50 5600 3150
rect 6000 3050 6250 3150
rect 6000 50 6100 3050
rect 6150 50 6250 3050
rect 6000 -50 6250 50
rect 6650 3050 6900 3150
rect 6650 50 6750 3050
rect 6800 50 6900 3050
rect 6650 -50 6900 50
rect 7300 -50 7350 3150
rect 7750 3050 8000 3150
rect 7750 50 7850 3050
rect 7900 50 8000 3050
rect 7750 -50 8000 50
rect 8650 3050 8900 3150
rect 8650 50 8750 3050
rect 8800 50 8900 3050
rect 8650 -50 8900 50
rect 9300 -50 9350 3150
rect 9750 3050 10000 3150
rect 9750 50 9850 3050
rect 9900 50 10000 3050
rect 9750 -50 10000 50
rect 10750 3050 11000 3150
rect 10750 50 10850 3050
rect 10900 50 11000 3050
rect 10750 -50 11000 50
rect 11400 -50 11450 3150
rect 11850 3050 12100 3150
rect 12350 3050 12600 3150
rect 11850 50 11950 3050
rect 12000 50 12100 3050
rect 12350 50 12450 3050
rect 12500 50 12600 3050
rect 11850 -50 12100 50
rect 12350 -50 12600 50
rect 13000 3050 13250 3150
rect 13000 50 13100 3050
rect 13150 50 13250 3050
rect 13000 -50 13250 50
<< ndiffc >>
rect -250 -3700 -200 -700
rect 400 -3700 450 -700
rect 900 -3700 950 -700
rect 1550 -3700 1600 -700
rect 2200 -3700 2250 -700
rect 2950 -3700 3000 -700
rect 3600 -3700 3650 -700
rect 4250 -3700 4300 -700
rect 5000 -3700 5050 -700
rect 6100 -3700 6150 -700
rect 6750 -3700 6800 -700
rect 7850 -3700 7900 -700
rect 8600 -3700 8650 -700
rect 9250 -3700 9300 -700
rect 9900 -3700 9950 -700
rect 10650 -3700 10700 -700
rect 11300 -3700 11350 -700
rect 11950 -3700 12000 -700
rect 12450 -3700 12500 -700
rect 13100 -3700 13150 -700
<< pdiffc >>
rect -250 50 -200 3050
rect 400 50 450 3050
rect 900 50 950 3050
rect 2000 50 2050 3050
rect 3000 50 3050 3050
rect 4100 50 4150 3050
rect 5000 50 5050 3050
rect 6100 50 6150 3050
rect 6750 50 6800 3050
rect 7850 50 7900 3050
rect 8750 50 8800 3050
rect 9850 50 9900 3050
rect 10850 50 10900 3050
rect 11950 50 12000 3050
rect 12450 50 12500 3050
rect 13100 50 13150 3050
<< psubdiff >>
rect -600 -700 -350 -600
rect -600 -3700 -500 -700
rect -450 -3700 -350 -700
rect -600 -3800 -350 -3700
rect 550 -700 800 -600
rect 550 -3700 650 -700
rect 700 -3700 800 -700
rect 550 -3800 800 -3700
rect 2600 -700 2850 -600
rect 2600 -3700 2700 -700
rect 2750 -3700 2850 -700
rect 2600 -3800 2850 -3700
rect 4650 -700 4900 -600
rect 4650 -3700 4750 -700
rect 4800 -3700 4900 -700
rect 4650 -3800 4900 -3700
rect 8000 -700 8250 -600
rect 8000 -3700 8100 -700
rect 8150 -3700 8250 -700
rect 8000 -3800 8250 -3700
rect 10050 -700 10300 -600
rect 10050 -3700 10150 -700
rect 10200 -3700 10300 -700
rect 10050 -3800 10300 -3700
rect 12100 -700 12350 -600
rect 12100 -3700 12200 -700
rect 12250 -3700 12350 -700
rect 12100 -3800 12350 -3700
rect 13250 -700 13500 -600
rect 13250 -3700 13350 -700
rect 13400 -3700 13500 -700
rect 13250 -3800 13500 -3700
<< nsubdiff >>
rect -600 3050 -350 3150
rect -600 50 -500 3050
rect -450 50 -350 3050
rect -600 -50 -350 50
rect 550 3050 800 3150
rect 550 50 650 3050
rect 700 50 800 3050
rect 550 -50 800 50
rect 2650 3050 2900 3150
rect 2650 50 2750 3050
rect 2800 50 2900 3050
rect 2650 -50 2900 50
rect 4650 3050 4900 3150
rect 4650 50 4750 3050
rect 4800 50 4900 3050
rect 4650 -50 4900 50
rect 8000 3050 8250 3150
rect 8000 50 8100 3050
rect 8150 50 8250 3050
rect 8000 -50 8250 50
rect 10000 3050 10250 3150
rect 10000 50 10100 3050
rect 10150 50 10250 3050
rect 10000 -50 10250 50
rect 12100 3050 12350 3150
rect 12100 50 12200 3050
rect 12250 50 12350 3050
rect 12100 -50 12350 50
rect 13250 3050 13500 3150
rect 13250 50 13350 3050
rect 13400 50 13500 3050
rect 13250 -50 13500 50
<< psubdiffcont >>
rect -500 -3700 -450 -700
rect 650 -3700 700 -700
rect 2700 -3700 2750 -700
rect 4750 -3700 4800 -700
rect 8100 -3700 8150 -700
rect 10150 -3700 10200 -700
rect 12200 -3700 12250 -700
rect 13350 -3700 13400 -700
<< nsubdiffcont >>
rect -500 50 -450 3050
rect 650 50 700 3050
rect 2750 50 2800 3050
rect 4750 50 4800 3050
rect 8100 50 8150 3050
rect 10100 50 10150 3050
rect 12200 50 12250 3050
rect 13350 50 13400 3050
<< poly >>
rect 1050 3200 11850 3300
rect -100 3150 300 3200
rect 1050 3150 1450 3200
rect 1500 3150 1900 3200
rect 3150 3150 3550 3200
rect 3600 3150 4000 3200
rect 5150 3150 5550 3200
rect 5600 3150 6000 3200
rect 6900 3150 7300 3200
rect 7350 3150 7750 3200
rect 8900 3150 9300 3200
rect 9350 3150 9750 3200
rect 11000 3150 11400 3200
rect 11450 3150 11850 3200
rect 12600 3150 13000 3200
rect -100 -100 300 -50
rect 1050 -100 1450 -50
rect 1500 -100 1900 -50
rect 3150 -100 3550 -50
rect 3600 -100 4000 -50
rect 5150 -100 5550 -50
rect 5600 -100 6000 -50
rect 6900 -100 7300 -50
rect 7350 -100 7750 -50
rect 8900 -100 9300 -50
rect 9350 -100 9750 -50
rect 11000 -100 11400 -50
rect 11450 -100 11850 -50
rect 12600 -100 13000 -50
rect -100 -150 50 -100
rect 12850 -150 13000 -100
rect -100 -200 -50 -150
rect 0 -200 50 -150
rect 2000 -200 2150 -150
rect 4100 -200 4250 -150
rect 8650 -200 8800 -150
rect 10750 -200 10900 -150
rect 12850 -200 12900 -150
rect 12950 -200 13000 -150
rect -100 -250 50 -200
rect 1350 -250 2050 -200
rect 2100 -250 2150 -200
rect 1350 -300 2150 -250
rect 3400 -250 4150 -200
rect 4200 -250 5400 -200
rect 3400 -300 5400 -250
rect 1350 -550 1450 -300
rect 3400 -550 3500 -300
rect 5300 -550 5400 -300
rect 7500 -250 8700 -200
rect 8750 -250 9500 -200
rect 7500 -300 9500 -250
rect 10750 -250 10800 -200
rect 10850 -250 11550 -200
rect 12850 -250 13000 -200
rect 10750 -300 11550 -250
rect 7500 -550 7600 -300
rect 9400 -550 9500 -300
rect 11450 -550 11550 -300
rect -100 -600 300 -550
rect 1050 -600 1450 -550
rect 1700 -600 2100 -550
rect 3100 -600 3500 -550
rect 3750 -600 4150 -550
rect 5150 -600 5550 -550
rect 5600 -600 6000 -550
rect 6900 -600 7300 -550
rect 7350 -600 7750 -550
rect 8750 -600 9150 -550
rect 9400 -600 9800 -550
rect 10800 -600 11200 -550
rect 11450 -600 11850 -550
rect 12600 -600 13000 -550
rect -100 -3850 300 -3800
rect 1050 -3850 1450 -3800
rect 1700 -3850 2100 -3800
rect 3100 -3850 3500 -3800
rect 3750 -3850 4150 -3800
rect 5150 -3850 5550 -3800
rect 5600 -3850 6000 -3800
rect 6900 -3850 7300 -3800
rect 7350 -3850 7750 -3800
rect 8750 -3850 9150 -3800
rect 9400 -3850 9800 -3800
rect 10800 -3850 11200 -3800
rect 11450 -3850 11850 -3800
rect 12600 -3850 13000 -3800
rect -100 -3900 50 -3850
rect -100 -3950 -50 -3900
rect 0 -3950 50 -3900
rect -100 -4000 50 -3950
rect 1150 -4000 1300 -3950
rect 1800 -4000 2000 -3850
rect 3850 -4000 4050 -3850
rect 5700 -4000 5900 -3850
rect 7000 -4000 7200 -3850
rect 8850 -4000 9050 -3850
rect 10900 -4000 11100 -3850
rect 12850 -3900 13000 -3850
rect 12850 -3950 12900 -3900
rect 12950 -3950 13000 -3900
rect 12850 -4000 13000 -3950
rect 1150 -4050 1200 -4000
rect 1250 -4050 11100 -4000
rect 1150 -4100 11100 -4050
rect 1150 -4200 3700 -4150
rect 1150 -4250 1200 -4200
rect 1250 -4250 3600 -4200
rect 3650 -4250 3700 -4200
rect 1150 -4300 1300 -4250
rect 3550 -4300 3700 -4250
<< polycont >>
rect -50 -200 0 -150
rect 12900 -200 12950 -150
rect 2050 -250 2100 -200
rect 4150 -250 4200 -200
rect 8700 -250 8750 -200
rect 10800 -250 10850 -200
rect -50 -3950 0 -3900
rect 12900 -3950 12950 -3900
rect 1200 -4050 1250 -4000
rect 1200 -4250 1250 -4200
rect 3600 -4250 3650 -4200
<< locali >>
rect -550 3100 -350 3150
rect 550 3100 800 3150
rect 2700 3100 2900 3150
rect 4700 3100 4900 3150
rect -550 3050 -150 3100
rect -550 50 -500 3050
rect -450 50 -250 3050
rect -200 50 -150 3050
rect -550 0 -150 50
rect 350 3050 1000 3100
rect 350 50 400 3050
rect 450 50 650 3050
rect 700 50 900 3050
rect 950 50 1000 3050
rect 350 0 1000 50
rect 1950 3050 2100 3100
rect 1950 50 2000 3050
rect 2050 50 2100 3050
rect 1950 0 2100 50
rect -550 -50 -350 0
rect -300 -100 -150 0
rect 550 -50 800 0
rect -300 -150 50 -100
rect -300 -200 -50 -150
rect 0 -200 50 -150
rect -300 -250 50 -200
rect 2000 -150 2100 0
rect 2700 3050 3100 3100
rect 2700 50 2750 3050
rect 2800 50 3000 3050
rect 3050 50 3100 3050
rect 2700 0 3100 50
rect 4050 3050 4200 3100
rect 4050 50 4100 3050
rect 4150 50 4200 3050
rect 4050 0 4200 50
rect 2700 -50 2900 0
rect 4100 -150 4200 0
rect 4700 3050 5100 3100
rect 4700 50 4750 3050
rect 4800 50 5000 3050
rect 5050 50 5100 3050
rect 4700 0 5100 50
rect 6050 3050 6200 3100
rect 6050 50 6100 3050
rect 6150 50 6200 3050
rect 4700 -50 4900 0
rect 2000 -200 2250 -150
rect 2000 -250 2050 -200
rect 2100 -250 2250 -200
rect 2000 -300 2250 -250
rect 4100 -200 4300 -150
rect 4100 -250 4150 -200
rect 4200 -250 4300 -200
rect 4100 -300 4300 -250
rect 2150 -650 2250 -300
rect 4200 -650 4300 -300
rect 6050 -300 6200 50
rect 6350 -300 6550 3400
rect 8000 3100 8200 3150
rect 10000 3100 10200 3150
rect 12100 3100 12350 3150
rect 13250 3100 13450 3150
rect 6700 3050 6850 3100
rect 6700 50 6750 3050
rect 6800 50 6850 3050
rect 6700 -300 6850 50
rect 7800 3050 8200 3100
rect 7800 50 7850 3050
rect 7900 50 8100 3050
rect 8150 50 8200 3050
rect 7800 0 8200 50
rect 8000 -50 8200 0
rect 8700 3050 8850 3100
rect 8700 50 8750 3050
rect 8800 50 8850 3050
rect 8700 0 8850 50
rect 9800 3050 10200 3100
rect 9800 50 9850 3050
rect 9900 50 10100 3050
rect 10150 50 10200 3050
rect 9800 0 10200 50
rect 8700 -150 8800 0
rect 10000 -50 10200 0
rect 10800 3050 10950 3100
rect 10800 50 10850 3050
rect 10900 50 10950 3050
rect 10800 0 10950 50
rect 11900 3050 12550 3100
rect 11900 50 11950 3050
rect 12000 50 12200 3050
rect 12250 50 12450 3050
rect 12500 50 12550 3050
rect 11900 0 12550 50
rect 13050 3050 13450 3100
rect 13050 50 13100 3050
rect 13150 50 13350 3050
rect 13400 50 13450 3050
rect 13050 0 13450 50
rect 10800 -150 10900 0
rect 12100 -50 12350 0
rect 13050 -100 13200 0
rect 13250 -50 13450 0
rect 6050 -400 6850 -300
rect -550 -700 -150 -650
rect -550 -3700 -500 -700
rect -450 -3700 -250 -700
rect -200 -3700 -150 -700
rect -550 -3750 -150 -3700
rect 350 -700 1000 -650
rect 350 -3700 400 -700
rect 450 -3700 650 -700
rect 700 -3700 900 -700
rect 950 -3700 1000 -700
rect 350 -3750 1000 -3700
rect 1500 -700 1650 -650
rect 1500 -3700 1550 -700
rect 1600 -3700 1650 -700
rect -300 -3850 -150 -3750
rect -300 -3900 50 -3850
rect -300 -3950 -50 -3900
rect 0 -3950 50 -3900
rect -300 -4000 50 -3950
rect 1150 -4000 1300 -3950
rect 250 -4050 1200 -4000
rect 1250 -4050 1300 -4000
rect -650 -4100 1300 -4050
rect -650 -4150 350 -4100
rect 1150 -4200 1300 -4150
rect -650 -4250 1200 -4200
rect 1250 -4250 1300 -4200
rect -650 -4300 1300 -4250
rect 1500 -4350 1650 -3700
rect 2150 -700 2300 -650
rect 2150 -3700 2200 -700
rect 2250 -3700 2300 -700
rect 2150 -3750 2300 -3700
rect 2650 -700 3050 -650
rect 2650 -3700 2700 -700
rect 2750 -3700 2950 -700
rect 3000 -3700 3050 -700
rect 2650 -3750 3050 -3700
rect 3550 -700 3700 -650
rect 3550 -3700 3600 -700
rect 3650 -3700 3700 -700
rect 3550 -4050 3700 -3700
rect 4200 -700 4350 -650
rect 4200 -3700 4250 -700
rect 4300 -3700 4350 -700
rect 4200 -3750 4350 -3700
rect 4700 -700 5100 -650
rect 4700 -3700 4750 -700
rect 4800 -3700 5000 -700
rect 5050 -3700 5100 -700
rect 4700 -3750 5100 -3700
rect 6050 -700 6200 -400
rect 6050 -3700 6100 -700
rect 6150 -3700 6200 -700
rect 6050 -3750 6200 -3700
rect 6700 -700 6850 -400
rect 8600 -200 8800 -150
rect 8600 -250 8700 -200
rect 8750 -250 8800 -200
rect 8600 -300 8800 -250
rect 10650 -200 10900 -150
rect 10650 -250 10800 -200
rect 10850 -250 10900 -200
rect 12850 -150 13200 -100
rect 12850 -200 12900 -150
rect 12950 -200 13200 -150
rect 12850 -250 13200 -200
rect 10650 -300 10900 -250
rect 8600 -650 8700 -300
rect 10650 -650 10750 -300
rect 6700 -3700 6750 -700
rect 6800 -3700 6850 -700
rect 6700 -3750 6850 -3700
rect 7800 -700 8200 -650
rect 7800 -3700 7850 -700
rect 7900 -3700 8100 -700
rect 8150 -3700 8200 -700
rect 7800 -3750 8200 -3700
rect 8550 -700 8700 -650
rect 8550 -3700 8600 -700
rect 8650 -3700 8700 -700
rect 8550 -3750 8700 -3700
rect 9200 -700 9350 -650
rect 9200 -3700 9250 -700
rect 9300 -3700 9350 -700
rect 9200 -4050 9350 -3700
rect 9850 -700 10250 -650
rect 9850 -3700 9900 -700
rect 9950 -3700 10150 -700
rect 10200 -3700 10250 -700
rect 9850 -3750 10250 -3700
rect 10600 -700 10750 -650
rect 10600 -3700 10650 -700
rect 10700 -3700 10750 -700
rect 10600 -3750 10750 -3700
rect 11250 -700 11400 -650
rect 11250 -3700 11300 -700
rect 11350 -3700 11400 -700
rect 3550 -4150 9350 -4050
rect 3550 -4200 3700 -4150
rect 3550 -4250 3600 -4200
rect 3650 -4250 3700 -4200
rect 3550 -4300 3700 -4250
rect 11250 -4350 11400 -3700
rect 11900 -700 12550 -650
rect 11900 -3700 11950 -700
rect 12000 -3700 12200 -700
rect 12250 -3700 12450 -700
rect 12500 -3700 12550 -700
rect 11900 -3750 12550 -3700
rect 13050 -700 13450 -650
rect 13050 -3700 13100 -700
rect 13150 -3700 13350 -700
rect 13400 -3700 13450 -700
rect 13050 -3750 13450 -3700
rect 13050 -3850 13200 -3750
rect 12850 -3900 13200 -3850
rect 12850 -3950 12900 -3900
rect 12950 -3950 13200 -3900
rect 12850 -4000 13200 -3950
rect -650 -4450 11400 -4350
<< viali >>
rect -500 50 -450 3050
rect 650 50 700 3050
rect 2750 50 2800 3050
rect 4750 50 4800 3050
rect 8100 50 8150 3050
rect 10100 50 10150 3050
rect 12200 50 12250 3050
rect 13350 50 13400 3050
rect -500 -3700 -450 -700
rect 650 -3700 700 -700
rect 2700 -3700 2750 -700
rect 4750 -3700 4800 -700
rect 8100 -3700 8150 -700
rect 10150 -3700 10200 -700
rect 12200 -3700 12250 -700
rect 13350 -3700 13400 -700
<< metal1 >>
rect -600 3050 -350 3150
rect -600 50 -500 3050
rect -450 50 -350 3050
rect -600 -50 -350 50
rect 550 3050 800 3150
rect 550 50 650 3050
rect 700 50 800 3050
rect 550 -50 800 50
rect 2650 3050 2900 3150
rect 2650 50 2750 3050
rect 2800 50 2900 3050
rect 2650 -50 2900 50
rect 4650 3050 4900 3150
rect 4650 50 4750 3050
rect 4800 50 4900 3050
rect 4650 -50 4900 50
rect 8000 3050 8250 3150
rect 8000 50 8100 3050
rect 8150 50 8250 3050
rect 8000 -50 8250 50
rect 10000 3050 10250 3150
rect 10000 50 10100 3050
rect 10150 50 10250 3050
rect 10000 -50 10250 50
rect 12100 3050 12350 3150
rect 12100 50 12200 3050
rect 12250 50 12350 3050
rect 12100 -50 12350 50
rect 13250 3050 13500 3150
rect 13250 50 13350 3050
rect 13400 50 13500 3050
rect 13250 -50 13500 50
rect -600 -200 13500 -50
rect -600 -700 -350 -650
rect -600 -3700 -500 -700
rect -450 -3700 -350 -700
rect -600 -3800 -350 -3700
rect 550 -700 800 -650
rect 550 -3700 650 -700
rect 700 -3700 800 -700
rect 550 -3800 800 -3700
rect 2600 -700 2850 -650
rect 2600 -3700 2700 -700
rect 2750 -3700 2850 -700
rect 2600 -3800 2850 -3700
rect 4650 -700 4900 -650
rect 4650 -3700 4750 -700
rect 4800 -3700 4900 -700
rect 4650 -3800 4900 -3700
rect 8000 -700 8250 -650
rect 8000 -3700 8100 -700
rect 8150 -3700 8250 -700
rect 8000 -3800 8250 -3700
rect 10050 -700 10300 -650
rect 10050 -3700 10150 -700
rect 10200 -3700 10300 -700
rect 10050 -3800 10300 -3700
rect 12100 -700 12350 -650
rect 12100 -3700 12200 -700
rect 12250 -3700 12350 -700
rect 12100 -3800 12350 -3700
rect 13250 -700 13500 -650
rect 13250 -3700 13350 -700
rect 13400 -3700 13500 -700
rect 13250 -3800 13500 -3700
rect -600 -3950 13500 -3800
<< labels >>
flabel locali -650 -4100 -650 -4100 0 FreeSans 240 0 0 0 VCN
port 0 nsew
flabel locali 6450 3400 6450 3400 0 FreeSans 240 0 0 0 i_fvf_out
port 3 nsew
flabel metal1 -600 -150 -600 -150 0 FreeSans 240 0 0 0 VDD
flabel metal1 -600 -3900 -600 -3900 0 FreeSans 240 0 0 0 GND
flabel locali -650 -4400 -650 -4400 0 FreeSans 240 0 0 0 i_dump
port 2 nsew
flabel locali -650 -4250 -650 -4250 0 FreeSans 240 0 0 0 i_out
port 1 nsew
<< end >>

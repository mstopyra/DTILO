magic
tech sky130A
magscale 1 2
timestamp 1702164466
<< error_p >>
rect -4700 -4400 -2360 -4350
rect -4700 -4509 -4699 -4460
rect -4700 -4510 -2360 -4509
rect -4700 -4620 -2360 -4570
rect -4700 -5040 -2360 -4990
<< nwell >>
rect -4830 -290 -1860 2600
rect -4870 -8070 -2230 -4070
<< nmos >>
rect -4660 -2940 -4560 -540
rect -4450 -2940 -4350 -540
rect -4300 -2940 -4200 -540
rect -4150 -2940 -4050 -540
rect -4000 -2940 -3900 -540
rect -3850 -2940 -3750 -540
rect -3640 -2940 -3540 -540
rect -3490 -2940 -3390 -540
rect -3340 -2940 -3240 -540
rect -3190 -2940 -3090 -540
rect -3040 -2940 -2940 -540
rect -2610 -2940 -2510 -540
rect -4730 -3370 -2330 -3270
rect -4730 -3800 -2330 -3700
rect -4670 -10750 -4570 -8350
rect -4460 -10750 -4360 -8350
rect -4250 -10750 -4150 -8350
rect -4040 -10750 -3940 -8350
rect -3830 -10750 -3730 -8350
rect -3620 -10750 -3520 -8350
rect -3190 -10750 -3090 -8350
rect -2980 -10750 -2880 -8350
rect -2770 -10750 -2670 -8350
rect -2560 -10750 -2460 -8350
rect -2350 -10750 -2250 -8350
rect -2140 -10750 -2040 -8350
<< pmos >>
rect -4660 -180 -4560 2220
rect -4450 -180 -4350 2220
rect -4240 -180 -4140 2220
rect -4030 -180 -3930 2220
rect -3820 -180 -3720 2220
rect -3610 -180 -3510 2220
rect -3180 -180 -3080 2220
rect -2970 -180 -2870 2220
rect -2760 -180 -2660 2220
rect -2550 -180 -2450 2220
rect -2340 -180 -2240 2220
rect -2130 -180 -2030 2220
rect -4730 -4320 -2330 -4220
rect -4730 -4750 -2330 -4650
rect -4730 -4960 -2330 -4860
rect -4730 -5170 -2330 -5070
rect -4670 -7990 -4570 -5590
rect -4460 -7990 -4360 -5590
rect -4310 -7990 -4210 -5590
rect -4160 -7990 -4060 -5590
rect -4010 -7990 -3910 -5590
rect -3860 -7990 -3760 -5590
rect -3650 -7990 -3550 -5590
rect -3500 -7990 -3400 -5590
rect -3350 -7990 -3250 -5590
rect -3200 -7990 -3100 -5590
rect -3050 -7990 -2950 -5590
rect -2620 -7990 -2520 -5590
<< ndiff >>
rect -4770 -570 -4660 -540
rect -4770 -2910 -4740 -570
rect -4690 -2910 -4660 -570
rect -4770 -2940 -4660 -2910
rect -4560 -570 -4450 -540
rect -4560 -2910 -4530 -570
rect -4480 -2910 -4450 -570
rect -4560 -2940 -4450 -2910
rect -4350 -2940 -4300 -540
rect -4200 -2940 -4150 -540
rect -4050 -2940 -4000 -540
rect -3900 -2940 -3850 -540
rect -3750 -570 -3640 -540
rect -3750 -2910 -3720 -570
rect -3670 -2910 -3640 -570
rect -3750 -2940 -3640 -2910
rect -3540 -2940 -3490 -540
rect -3390 -2940 -3340 -540
rect -3240 -2940 -3190 -540
rect -3090 -2940 -3040 -540
rect -2940 -570 -2830 -540
rect -2720 -570 -2610 -540
rect -2940 -2910 -2910 -570
rect -2860 -2910 -2830 -570
rect -2720 -2910 -2690 -570
rect -2640 -2910 -2610 -570
rect -2940 -2940 -2830 -2910
rect -2720 -2940 -2610 -2910
rect -2510 -570 -2400 -540
rect -2510 -2910 -2480 -570
rect -2430 -2910 -2400 -570
rect -2510 -2940 -2400 -2910
rect -4730 -3190 -2330 -3160
rect -4730 -3240 -4700 -3190
rect -2360 -3240 -2330 -3190
rect -4730 -3270 -2330 -3240
rect -4730 -3400 -2330 -3370
rect -4730 -3450 -4700 -3400
rect -2360 -3450 -2330 -3400
rect -4730 -3480 -2330 -3450
rect -4730 -3620 -2330 -3590
rect -4730 -3670 -4700 -3620
rect -2360 -3670 -2330 -3620
rect -4730 -3700 -2330 -3670
rect -4730 -3830 -2330 -3800
rect -4730 -3880 -4700 -3830
rect -2360 -3880 -2330 -3830
rect -4730 -3910 -2330 -3880
rect -4780 -8380 -4670 -8350
rect -4780 -10720 -4750 -8380
rect -4700 -10720 -4670 -8380
rect -4780 -10750 -4670 -10720
rect -4570 -8380 -4460 -8350
rect -4570 -10720 -4540 -8380
rect -4490 -10720 -4460 -8380
rect -4570 -10750 -4460 -10720
rect -4360 -8380 -4250 -8350
rect -4360 -10720 -4330 -8380
rect -4280 -10720 -4250 -8380
rect -4360 -10750 -4250 -10720
rect -4150 -8380 -4040 -8350
rect -4150 -10720 -4120 -8380
rect -4070 -10720 -4040 -8380
rect -4150 -10750 -4040 -10720
rect -3940 -8380 -3830 -8350
rect -3940 -10720 -3910 -8380
rect -3860 -10720 -3830 -8380
rect -3940 -10750 -3830 -10720
rect -3730 -8380 -3620 -8350
rect -3730 -10720 -3700 -8380
rect -3650 -10720 -3620 -8380
rect -3730 -10750 -3620 -10720
rect -3520 -8380 -3410 -8350
rect -3300 -8380 -3190 -8350
rect -3520 -10720 -3490 -8380
rect -3440 -10720 -3410 -8380
rect -3300 -10720 -3270 -8380
rect -3220 -10720 -3190 -8380
rect -3520 -10750 -3410 -10720
rect -3300 -10750 -3190 -10720
rect -3090 -8380 -2980 -8350
rect -3090 -10720 -3060 -8380
rect -3010 -10720 -2980 -8380
rect -3090 -10750 -2980 -10720
rect -2880 -8380 -2770 -8350
rect -2880 -10720 -2850 -8380
rect -2800 -10720 -2770 -8380
rect -2880 -10750 -2770 -10720
rect -2670 -8380 -2560 -8350
rect -2670 -10720 -2640 -8380
rect -2590 -10720 -2560 -8380
rect -2670 -10750 -2560 -10720
rect -2460 -8380 -2350 -8350
rect -2460 -10720 -2430 -8380
rect -2380 -10720 -2350 -8380
rect -2460 -10750 -2350 -10720
rect -2250 -8380 -2140 -8350
rect -2250 -10720 -2220 -8380
rect -2170 -10720 -2140 -8380
rect -2250 -10750 -2140 -10720
rect -2040 -8380 -1930 -8350
rect -2040 -10720 -2010 -8380
rect -1960 -10720 -1930 -8380
rect -2040 -10750 -1930 -10720
<< pdiff >>
rect -4770 2190 -4660 2220
rect -4770 -150 -4740 2190
rect -4690 -150 -4660 2190
rect -4770 -180 -4660 -150
rect -4560 2190 -4450 2220
rect -4560 -150 -4530 2190
rect -4480 -150 -4450 2190
rect -4560 -180 -4450 -150
rect -4350 2190 -4240 2220
rect -4350 -150 -4320 2190
rect -4270 -150 -4240 2190
rect -4350 -180 -4240 -150
rect -4140 2190 -4030 2220
rect -4140 -150 -4110 2190
rect -4060 -150 -4030 2190
rect -4140 -180 -4030 -150
rect -3930 2190 -3820 2220
rect -3930 -150 -3900 2190
rect -3850 -150 -3820 2190
rect -3930 -180 -3820 -150
rect -3720 2190 -3610 2220
rect -3720 -150 -3690 2190
rect -3640 -150 -3610 2190
rect -3720 -180 -3610 -150
rect -3510 2190 -3400 2220
rect -3290 2190 -3180 2220
rect -3510 -150 -3480 2190
rect -3430 -150 -3400 2190
rect -3290 -150 -3260 2190
rect -3210 -150 -3180 2190
rect -3510 -180 -3400 -150
rect -3290 -180 -3180 -150
rect -3080 2190 -2970 2220
rect -3080 -150 -3050 2190
rect -3000 -150 -2970 2190
rect -3080 -180 -2970 -150
rect -2870 2190 -2760 2220
rect -2870 -150 -2840 2190
rect -2790 -150 -2760 2190
rect -2870 -180 -2760 -150
rect -2660 2190 -2550 2220
rect -2660 -150 -2630 2190
rect -2580 -150 -2550 2190
rect -2660 -180 -2550 -150
rect -2450 2190 -2340 2220
rect -2450 -150 -2420 2190
rect -2370 -150 -2340 2190
rect -2450 -180 -2340 -150
rect -2240 2190 -2130 2220
rect -2240 -150 -2210 2190
rect -2160 -150 -2130 2190
rect -2240 -180 -2130 -150
rect -2030 2190 -1920 2220
rect -2030 -150 -2000 2190
rect -1950 -150 -1920 2190
rect -2030 -180 -1920 -150
rect -4730 -4140 -2330 -4110
rect -4730 -4190 -4700 -4140
rect -2360 -4190 -2330 -4140
rect -4730 -4220 -2330 -4190
rect -4730 -4350 -2330 -4320
rect -4730 -4400 -4700 -4350
rect -2360 -4400 -2330 -4350
rect -4730 -4430 -2330 -4400
rect -4730 -4570 -2330 -4540
rect -4730 -4620 -4700 -4570
rect -2360 -4620 -2330 -4570
rect -4730 -4650 -2330 -4620
rect -4730 -4780 -2330 -4750
rect -4730 -4830 -4700 -4780
rect -2360 -4830 -2330 -4780
rect -4730 -4860 -2330 -4830
rect -4730 -4990 -2330 -4960
rect -4730 -5040 -4700 -4990
rect -2360 -5040 -2330 -4990
rect -4730 -5070 -2330 -5040
rect -4730 -5200 -2330 -5170
rect -4730 -5250 -4700 -5200
rect -2360 -5250 -2330 -5200
rect -4730 -5280 -2330 -5250
rect -4780 -5620 -4670 -5590
rect -4780 -7960 -4750 -5620
rect -4700 -7960 -4670 -5620
rect -4780 -7990 -4670 -7960
rect -4570 -5620 -4460 -5590
rect -4570 -7960 -4540 -5620
rect -4490 -7960 -4460 -5620
rect -4570 -7990 -4460 -7960
rect -4360 -7990 -4310 -5590
rect -4210 -7990 -4160 -5590
rect -4060 -7990 -4010 -5590
rect -3910 -7990 -3860 -5590
rect -3760 -5620 -3650 -5590
rect -3760 -7960 -3730 -5620
rect -3680 -7960 -3650 -5620
rect -3760 -7990 -3650 -7960
rect -3550 -7990 -3500 -5590
rect -3400 -7990 -3350 -5590
rect -3250 -7990 -3200 -5590
rect -3100 -7990 -3050 -5590
rect -2950 -5620 -2840 -5590
rect -2730 -5620 -2620 -5590
rect -2950 -7960 -2920 -5620
rect -2870 -7960 -2840 -5620
rect -2730 -7960 -2700 -5620
rect -2650 -7960 -2620 -5620
rect -2950 -7990 -2840 -7960
rect -2730 -7990 -2620 -7960
rect -2520 -5620 -2410 -5590
rect -2520 -7960 -2490 -5620
rect -2440 -7960 -2410 -5620
rect -2520 -7990 -2410 -7960
<< ndiffc >>
rect -4740 -2910 -4690 -570
rect -4530 -2910 -4480 -570
rect -3720 -2910 -3670 -570
rect -2910 -2910 -2860 -570
rect -2690 -2910 -2640 -570
rect -2480 -2910 -2430 -570
rect -4700 -3240 -2360 -3190
rect -4700 -3450 -2360 -3400
rect -4700 -3670 -2360 -3620
rect -4700 -3880 -2360 -3830
rect -4750 -10720 -4700 -8380
rect -4540 -10720 -4490 -8380
rect -4330 -10720 -4280 -8380
rect -4120 -10720 -4070 -8380
rect -3910 -10720 -3860 -8380
rect -3700 -10720 -3650 -8380
rect -3490 -10720 -3440 -8380
rect -3270 -10720 -3220 -8380
rect -3060 -10720 -3010 -8380
rect -2850 -10720 -2800 -8380
rect -2640 -10720 -2590 -8380
rect -2430 -10720 -2380 -8380
rect -2220 -10720 -2170 -8380
rect -2010 -10720 -1960 -8380
<< pdiffc >>
rect -4740 -150 -4690 2190
rect -4530 -150 -4480 2190
rect -4320 -150 -4270 2190
rect -4110 -150 -4060 2190
rect -3900 -150 -3850 2190
rect -3690 -150 -3640 2190
rect -3480 -150 -3430 2190
rect -3260 -150 -3210 2190
rect -3050 -150 -3000 2190
rect -2840 -150 -2790 2190
rect -2630 -150 -2580 2190
rect -2420 -150 -2370 2190
rect -2210 -150 -2160 2190
rect -2000 -150 -1950 2190
rect -4700 -4190 -2360 -4140
rect -4700 -4400 -2360 -4350
rect -4700 -4620 -2360 -4570
rect -4700 -4830 -2360 -4780
rect -4700 -5040 -2360 -4990
rect -4700 -5250 -2360 -5200
rect -4750 -7960 -4700 -5620
rect -4540 -7960 -4490 -5620
rect -3730 -7960 -3680 -5620
rect -2920 -7960 -2870 -5620
rect -2700 -7960 -2650 -5620
rect -2490 -7960 -2440 -5620
<< psubdiff >>
rect -2830 -570 -2720 -540
rect -2830 -2910 -2800 -570
rect -2750 -2910 -2720 -570
rect -2830 -2940 -2720 -2910
rect -4730 -3510 -2330 -3480
rect -4730 -3560 -4700 -3510
rect -2360 -3560 -2330 -3510
rect -4730 -3590 -2330 -3560
rect -3410 -8380 -3300 -8350
rect -3410 -10720 -3380 -8380
rect -3330 -10720 -3300 -8380
rect -3410 -10750 -3300 -10720
<< nsubdiff >>
rect -3400 2190 -3290 2220
rect -3400 -150 -3370 2190
rect -3320 -150 -3290 2190
rect -3400 -180 -3290 -150
rect -4730 -4460 -2330 -4430
rect -4730 -4510 -4700 -4460
rect -2360 -4510 -2330 -4460
rect -4730 -4540 -2330 -4510
rect -2840 -5620 -2730 -5590
rect -2840 -7960 -2810 -5620
rect -2760 -7960 -2730 -5620
rect -2840 -7990 -2730 -7960
<< psubdiffcont >>
rect -2800 -2910 -2750 -570
rect -4700 -3560 -2360 -3510
rect -3380 -10720 -3330 -8380
<< nsubdiffcont >>
rect -3370 -150 -3320 2190
rect -4700 -4510 -2360 -4460
rect -2810 -7960 -2760 -5620
<< poly >>
rect -4660 2220 -4560 2250
rect -4450 2220 -4350 2250
rect -4240 2220 -4140 2250
rect -4030 2220 -3930 2250
rect -3820 2220 -3720 2250
rect -3610 2220 -3510 2250
rect -3180 2220 -3080 2250
rect -2970 2220 -2870 2250
rect -2760 2220 -2660 2250
rect -2550 2220 -2450 2250
rect -2340 2220 -2240 2250
rect -2130 2220 -2030 2250
rect -4660 -320 -4560 -180
rect -4450 -210 -4350 -180
rect -4240 -210 -4140 -180
rect -4030 -210 -3930 -180
rect -3820 -210 -3720 -180
rect -3610 -210 -3510 -180
rect -3180 -210 -3080 -180
rect -2970 -210 -2870 -180
rect -2760 -210 -2660 -180
rect -2550 -210 -2450 -180
rect -2340 -210 -2240 -180
rect -4450 -230 -2240 -210
rect -4450 -290 -4330 -230
rect -4260 -290 -4120 -230
rect -4050 -290 -3910 -230
rect -3840 -290 -3490 -230
rect -3420 -290 -2850 -230
rect -2780 -290 -2640 -230
rect -2570 -290 -2430 -230
rect -2360 -290 -2240 -230
rect -4450 -310 -2240 -290
rect -4760 -340 -4560 -320
rect -4760 -400 -4740 -340
rect -4680 -400 -4560 -340
rect -2130 -360 -2030 -180
rect -4760 -420 -4560 -400
rect -2250 -380 -2030 -360
rect -2250 -440 -2230 -380
rect -2170 -440 -2030 -380
rect -2250 -460 -2030 -440
rect -4660 -540 -4560 -510
rect -4450 -540 -4350 -510
rect -4300 -540 -4200 -510
rect -4150 -540 -4050 -510
rect -4000 -540 -3900 -510
rect -3850 -540 -3750 -510
rect -3640 -540 -3540 -510
rect -3490 -540 -3390 -510
rect -3340 -540 -3240 -510
rect -3190 -540 -3090 -510
rect -3040 -540 -2940 -510
rect -2610 -540 -2510 -510
rect -4660 -2970 -4560 -2940
rect -4450 -2970 -4350 -2940
rect -4300 -2970 -4200 -2940
rect -4150 -2970 -4050 -2940
rect -4000 -2970 -3900 -2940
rect -3850 -2970 -3750 -2940
rect -3640 -2970 -3540 -2940
rect -3490 -2970 -3390 -2940
rect -3340 -2970 -3240 -2940
rect -3190 -2970 -3090 -2940
rect -3040 -2970 -2940 -2940
rect -2610 -2970 -2510 -2940
rect -4850 -3070 -2510 -2970
rect -4850 -3270 -4750 -3070
rect -4850 -3370 -4730 -3270
rect -2330 -3290 -2200 -3270
rect -2330 -3350 -2280 -3290
rect -2220 -3350 -2200 -3290
rect -2330 -3370 -2200 -3350
rect -4760 -3800 -4730 -3700
rect -2330 -3720 -2200 -3700
rect -2330 -3780 -2280 -3720
rect -2220 -3780 -2200 -3720
rect -2330 -3800 -2200 -3780
rect -4870 -4320 -4730 -4220
rect -2330 -4320 -2300 -4220
rect -4870 -4650 -4760 -4320
rect -4870 -4750 -4730 -4650
rect -2330 -4750 -2300 -4650
rect -4870 -4860 -4760 -4750
rect -4870 -4960 -4730 -4860
rect -2330 -4960 -2300 -4860
rect -4870 -5070 -4760 -4960
rect -4870 -5170 -4730 -5070
rect -2330 -5090 -2200 -5070
rect -2330 -5150 -2280 -5090
rect -2220 -5150 -2200 -5090
rect -2330 -5170 -2200 -5150
rect -4870 -5360 -4760 -5170
rect -4870 -5380 -4570 -5360
rect -4870 -5440 -4650 -5380
rect -4590 -5440 -4570 -5380
rect -4870 -5450 -4570 -5440
rect -4670 -5460 -4570 -5450
rect -4670 -5560 -2520 -5460
rect -4670 -5590 -4570 -5560
rect -4460 -5590 -4360 -5560
rect -4310 -5590 -4210 -5560
rect -4160 -5590 -4060 -5560
rect -4010 -5590 -3910 -5560
rect -3860 -5590 -3760 -5560
rect -3650 -5590 -3550 -5560
rect -3500 -5590 -3400 -5560
rect -3350 -5590 -3250 -5560
rect -3200 -5590 -3100 -5560
rect -3050 -5590 -2950 -5560
rect -2620 -5590 -2520 -5560
rect -4670 -8020 -4570 -7990
rect -4460 -8020 -4360 -7990
rect -4310 -8020 -4210 -7990
rect -4160 -8020 -4060 -7990
rect -4010 -8020 -3910 -7990
rect -3860 -8020 -3760 -7990
rect -3650 -8020 -3550 -7990
rect -3500 -8020 -3400 -7990
rect -3350 -8020 -3250 -7990
rect -3200 -8020 -3100 -7990
rect -3050 -8020 -2950 -7990
rect -2620 -8020 -2520 -7990
rect -2260 -8090 -2040 -8070
rect -4770 -8130 -4570 -8110
rect -4770 -8190 -4750 -8130
rect -4690 -8190 -4570 -8130
rect -2260 -8150 -2240 -8090
rect -2180 -8150 -2040 -8090
rect -2260 -8170 -2040 -8150
rect -4770 -8210 -4570 -8190
rect -4670 -8350 -4570 -8210
rect -4460 -8240 -2250 -8220
rect -4460 -8300 -4340 -8240
rect -4270 -8300 -4130 -8240
rect -4060 -8300 -3920 -8240
rect -3850 -8300 -3500 -8240
rect -3430 -8300 -2860 -8240
rect -2790 -8300 -2650 -8240
rect -2580 -8300 -2440 -8240
rect -2370 -8300 -2250 -8240
rect -4460 -8320 -2250 -8300
rect -4460 -8350 -4360 -8320
rect -4250 -8350 -4150 -8320
rect -4040 -8350 -3940 -8320
rect -3830 -8350 -3730 -8320
rect -3620 -8350 -3520 -8320
rect -3190 -8350 -3090 -8320
rect -2980 -8350 -2880 -8320
rect -2770 -8350 -2670 -8320
rect -2560 -8350 -2460 -8320
rect -2350 -8350 -2250 -8320
rect -2140 -8350 -2040 -8170
rect -4670 -10780 -4570 -10750
rect -4460 -10780 -4360 -10750
rect -4250 -10780 -4150 -10750
rect -4040 -10780 -3940 -10750
rect -3830 -10780 -3730 -10750
rect -3620 -10780 -3520 -10750
rect -3190 -10780 -3090 -10750
rect -2980 -10780 -2880 -10750
rect -2770 -10780 -2670 -10750
rect -2560 -10780 -2460 -10750
rect -2350 -10780 -2250 -10750
rect -2140 -10780 -2040 -10750
<< polycont >>
rect -4330 -290 -4260 -230
rect -4120 -290 -4050 -230
rect -3910 -290 -3840 -230
rect -3490 -290 -3420 -230
rect -2850 -290 -2780 -230
rect -2640 -290 -2570 -230
rect -2430 -290 -2360 -230
rect -4740 -400 -4680 -340
rect -2230 -440 -2170 -380
rect -2280 -3350 -2220 -3290
rect -2280 -3780 -2220 -3720
rect -2280 -5150 -2220 -5090
rect -4650 -5440 -4590 -5380
rect -4750 -8190 -4690 -8130
rect -2240 -8150 -2180 -8090
rect -4340 -8300 -4270 -8240
rect -4130 -8300 -4060 -8240
rect -3920 -8300 -3850 -8240
rect -3500 -8300 -3430 -8240
rect -2860 -8300 -2790 -8240
rect -2650 -8300 -2580 -8240
rect -2440 -8300 -2370 -8240
<< locali >>
rect -4940 2460 -1930 2550
rect -4940 2410 -4670 2460
rect -4760 2190 -4670 2410
rect -4760 -150 -4740 2190
rect -4690 -150 -4670 2190
rect -4760 -320 -4670 -150
rect -4550 2300 -2140 2390
rect -4550 2190 -4460 2300
rect -4550 -150 -4530 2190
rect -4480 -150 -4460 2190
rect -4550 -170 -4460 -150
rect -4340 2190 -4250 2210
rect -4340 -150 -4320 2190
rect -4270 -150 -4250 2190
rect -4340 -210 -4250 -150
rect -4130 2190 -4040 2210
rect -4130 -150 -4110 2190
rect -4060 -150 -4040 2190
rect -4130 -210 -4040 -150
rect -3920 2190 -3830 2210
rect -3920 -150 -3900 2190
rect -3850 -150 -3830 2190
rect -3920 -210 -3830 -150
rect -3710 2190 -3620 2300
rect -3710 -150 -3690 2190
rect -3640 -150 -3620 2190
rect -3710 -170 -3620 -150
rect -3500 2190 -3190 2210
rect -3500 -150 -3480 2190
rect -3430 -150 -3370 2190
rect -3320 -150 -3260 2190
rect -3210 -150 -3190 2190
rect -3500 -170 -3190 -150
rect -3070 2190 -2980 2300
rect -3070 -150 -3050 2190
rect -3000 -150 -2980 2190
rect -3070 -170 -2980 -150
rect -2860 2190 -2770 2210
rect -2860 -150 -2840 2190
rect -2790 -150 -2770 2190
rect -2860 -210 -2770 -150
rect -2650 2190 -2560 2210
rect -2650 -150 -2630 2190
rect -2580 -150 -2560 2190
rect -2650 -210 -2560 -150
rect -2440 2190 -2350 2210
rect -2440 -150 -2420 2190
rect -2370 -150 -2350 2190
rect -2440 -210 -2350 -150
rect -2230 2190 -2140 2300
rect -2230 -150 -2210 2190
rect -2160 -150 -2140 2190
rect -2230 -170 -2140 -150
rect -2020 2190 -1930 2460
rect -2020 -150 -2000 2190
rect -1950 -150 -1930 2190
rect -4350 -230 -4240 -210
rect -4350 -290 -4330 -230
rect -4260 -290 -4240 -230
rect -4350 -310 -4240 -290
rect -4140 -230 -4030 -210
rect -4140 -290 -4120 -230
rect -4050 -290 -4030 -230
rect -4140 -310 -4030 -290
rect -3930 -230 -3820 -210
rect -3930 -290 -3910 -230
rect -3840 -290 -3820 -230
rect -3930 -310 -3820 -290
rect -3510 -230 -3400 -210
rect -3510 -290 -3490 -230
rect -3420 -290 -3400 -230
rect -3510 -310 -3400 -290
rect -2870 -230 -2760 -210
rect -2870 -290 -2850 -230
rect -2780 -290 -2760 -230
rect -2870 -310 -2760 -290
rect -2660 -230 -2550 -210
rect -2660 -290 -2640 -230
rect -2570 -290 -2550 -230
rect -2660 -310 -2550 -290
rect -2450 -230 -2340 -210
rect -2450 -290 -2430 -230
rect -2360 -290 -2340 -230
rect -2450 -310 -2340 -290
rect -4760 -340 -4660 -320
rect -4760 -400 -4740 -340
rect -4680 -400 -4660 -340
rect -3510 -350 -3420 -310
rect -4760 -420 -4660 -400
rect -4760 -570 -4670 -420
rect -3740 -440 -3420 -350
rect -2250 -370 -2150 -360
rect -2020 -370 -1930 -150
rect -2500 -380 -1930 -370
rect -2500 -440 -2230 -380
rect -2170 -440 -1930 -380
rect -4760 -2910 -4740 -570
rect -4690 -2910 -4670 -570
rect -4760 -2930 -4670 -2910
rect -4550 -570 -4460 -550
rect -4550 -2910 -4530 -570
rect -4480 -2910 -4460 -570
rect -4550 -2930 -4460 -2910
rect -3740 -570 -3650 -440
rect -2500 -460 -1930 -440
rect -3740 -2910 -3720 -570
rect -3670 -2910 -3650 -570
rect -3740 -2930 -3650 -2910
rect -2930 -570 -2620 -550
rect -2930 -2910 -2910 -570
rect -2860 -2910 -2800 -570
rect -2750 -2910 -2690 -570
rect -2640 -2910 -2620 -570
rect -2930 -2930 -2620 -2910
rect -2500 -570 -2410 -460
rect -2500 -2910 -2480 -570
rect -2430 -2910 -2410 -570
rect -2500 -2930 -2410 -2910
rect -4930 -3170 -4840 -3020
rect -4930 -3190 -2200 -3170
rect -4930 -3240 -4700 -3190
rect -2360 -3240 -2200 -3190
rect -4930 -3260 -2200 -3240
rect -4930 -3810 -4840 -3260
rect -2300 -3290 -2200 -3260
rect -2300 -3350 -2280 -3290
rect -2220 -3350 -2200 -3290
rect -2300 -3370 -2200 -3350
rect -4720 -3400 -2340 -3380
rect -4720 -3450 -4700 -3400
rect -2360 -3450 -2340 -3400
rect -4720 -3510 -2340 -3450
rect -4720 -3560 -4700 -3510
rect -2360 -3560 -2340 -3510
rect -4720 -3620 -2340 -3560
rect -4720 -3670 -4700 -3620
rect -2360 -3670 -2340 -3620
rect -4720 -3690 -2340 -3670
rect -2300 -3720 -2200 -3700
rect -2300 -3780 -2280 -3720
rect -2220 -3780 -2200 -3720
rect -2300 -3810 -2200 -3780
rect -4930 -3830 -2200 -3810
rect -4930 -3880 -4700 -3830
rect -2360 -3880 -2200 -3830
rect -4930 -3900 -2200 -3880
rect -4930 -4760 -4840 -3900
rect -4720 -4140 -2340 -4120
rect -4720 -4190 -4700 -4140
rect -2360 -4190 -2340 -4140
rect -4720 -4210 -2340 -4190
rect -4720 -4350 -2340 -4330
rect -4720 -4400 -4700 -4350
rect -2360 -4400 -2340 -4350
rect -4720 -4460 -2340 -4400
rect -4720 -4510 -4700 -4460
rect -2360 -4510 -2340 -4460
rect -4720 -4570 -2340 -4510
rect -4720 -4620 -4700 -4570
rect -2360 -4620 -2340 -4570
rect -4720 -4640 -2340 -4620
rect -4930 -4780 -2330 -4760
rect -4930 -4830 -4700 -4780
rect -2360 -4830 -2330 -4780
rect -4930 -4850 -2330 -4830
rect -4720 -4990 -2340 -4970
rect -4720 -5040 -4700 -4990
rect -2360 -5040 -2340 -4990
rect -4720 -5060 -2340 -5040
rect -2300 -5090 -2200 -5070
rect -2300 -5150 -2280 -5090
rect -2220 -5150 -2200 -5090
rect -2300 -5180 -2200 -5150
rect -4720 -5200 -2200 -5180
rect -4720 -5250 -4700 -5200
rect -2360 -5250 -2200 -5200
rect -4720 -5270 -2200 -5250
rect -4940 -5380 -4570 -5360
rect -4940 -5440 -4650 -5380
rect -4590 -5440 -4570 -5380
rect -4940 -5450 -4570 -5440
rect -4670 -5460 -4570 -5450
rect -4770 -5620 -4680 -5600
rect -4770 -7960 -4750 -5620
rect -4700 -7960 -4680 -5620
rect -4770 -8110 -4680 -7960
rect -4560 -5620 -4470 -5600
rect -4560 -7960 -4540 -5620
rect -4490 -7960 -4470 -5620
rect -4560 -7980 -4470 -7960
rect -3750 -5620 -3660 -5600
rect -3750 -7960 -3730 -5620
rect -3680 -7960 -3660 -5620
rect -3750 -8090 -3660 -7960
rect -2940 -5620 -2630 -5600
rect -2940 -7960 -2920 -5620
rect -2870 -7960 -2810 -5620
rect -2760 -7960 -2700 -5620
rect -2650 -7960 -2630 -5620
rect -2940 -7980 -2630 -7960
rect -2510 -5620 -2420 -5600
rect -2510 -7960 -2490 -5620
rect -2440 -7960 -2420 -5620
rect -2510 -8070 -2420 -7960
rect -2510 -8090 -1940 -8070
rect -4770 -8130 -4670 -8110
rect -4770 -8190 -4750 -8130
rect -4690 -8190 -4670 -8130
rect -3750 -8180 -3430 -8090
rect -2510 -8150 -2240 -8090
rect -2180 -8150 -1940 -8090
rect -2510 -8160 -1940 -8150
rect -2260 -8170 -2160 -8160
rect -4770 -8210 -4670 -8190
rect -4770 -8380 -4680 -8210
rect -3520 -8220 -3430 -8180
rect -4360 -8240 -4250 -8220
rect -4360 -8300 -4340 -8240
rect -4270 -8300 -4250 -8240
rect -4360 -8320 -4250 -8300
rect -4150 -8240 -4040 -8220
rect -4150 -8300 -4130 -8240
rect -4060 -8300 -4040 -8240
rect -4150 -8320 -4040 -8300
rect -3940 -8240 -3830 -8220
rect -3940 -8300 -3920 -8240
rect -3850 -8300 -3830 -8240
rect -3940 -8320 -3830 -8300
rect -3520 -8240 -3410 -8220
rect -3520 -8300 -3500 -8240
rect -3430 -8300 -3410 -8240
rect -3520 -8320 -3410 -8300
rect -2880 -8240 -2770 -8220
rect -2880 -8300 -2860 -8240
rect -2790 -8300 -2770 -8240
rect -2880 -8320 -2770 -8300
rect -2670 -8240 -2560 -8220
rect -2670 -8300 -2650 -8240
rect -2580 -8300 -2560 -8240
rect -2670 -8320 -2560 -8300
rect -2460 -8240 -2350 -8220
rect -2460 -8300 -2440 -8240
rect -2370 -8300 -2350 -8240
rect -2460 -8320 -2350 -8300
rect -4770 -10720 -4750 -8380
rect -4700 -10720 -4680 -8380
rect -4770 -10930 -4680 -10720
rect -4560 -8380 -4470 -8360
rect -4560 -10720 -4540 -8380
rect -4490 -10720 -4470 -8380
rect -4560 -10830 -4470 -10720
rect -4350 -8380 -4260 -8320
rect -4350 -10720 -4330 -8380
rect -4280 -10720 -4260 -8380
rect -4350 -10740 -4260 -10720
rect -4140 -8380 -4050 -8320
rect -4140 -10720 -4120 -8380
rect -4070 -10720 -4050 -8380
rect -4140 -10740 -4050 -10720
rect -3930 -8380 -3840 -8320
rect -3930 -10720 -3910 -8380
rect -3860 -10720 -3840 -8380
rect -3930 -10740 -3840 -10720
rect -3720 -8380 -3630 -8360
rect -3720 -10720 -3700 -8380
rect -3650 -10720 -3630 -8380
rect -3720 -10830 -3630 -10720
rect -3510 -8380 -3200 -8360
rect -3510 -10720 -3490 -8380
rect -3440 -10720 -3380 -8380
rect -3330 -10720 -3270 -8380
rect -3220 -10720 -3200 -8380
rect -3510 -10740 -3200 -10720
rect -3080 -8380 -2990 -8360
rect -3080 -10720 -3060 -8380
rect -3010 -10720 -2990 -8380
rect -3080 -10830 -2990 -10720
rect -2870 -8380 -2780 -8320
rect -2870 -10720 -2850 -8380
rect -2800 -10720 -2780 -8380
rect -2870 -10740 -2780 -10720
rect -2660 -8380 -2570 -8320
rect -2660 -10720 -2640 -8380
rect -2590 -10720 -2570 -8380
rect -2660 -10740 -2570 -10720
rect -2450 -8380 -2360 -8320
rect -2450 -10720 -2430 -8380
rect -2380 -10720 -2360 -8380
rect -2450 -10740 -2360 -10720
rect -2240 -8380 -2150 -8360
rect -2240 -10720 -2220 -8380
rect -2170 -10720 -2150 -8380
rect -2240 -10830 -2150 -10720
rect -4560 -10920 -2150 -10830
rect -2030 -8380 -1940 -8160
rect -2030 -10720 -2010 -8380
rect -1960 -10720 -1940 -8380
rect -4940 -10990 -4680 -10930
rect -2030 -10990 -1940 -10720
rect -4940 -11080 -1940 -10990
<< viali >>
rect -3480 600 -3430 1810
rect -3370 600 -3320 1810
rect -3260 600 -3210 1810
rect -4530 -2250 -4480 -880
rect -2910 -2250 -2860 -880
rect -2800 -2250 -2750 -880
rect -2690 -2250 -2640 -880
rect -4700 -3450 -2360 -3400
rect -4700 -3560 -2360 -3510
rect -4700 -3670 -2360 -3620
rect -4700 -4400 -2360 -4350
rect -4700 -4510 -2360 -4460
rect -4700 -4620 -2360 -4570
rect -4700 -5040 -2360 -4990
rect -4540 -7460 -4490 -6080
rect -2920 -7460 -2870 -6080
rect -2810 -7460 -2760 -6080
rect -2700 -7460 -2650 -6080
rect -3490 -10180 -3440 -8950
rect -3380 -10180 -3330 -8950
rect -3270 -10180 -3220 -8950
<< metal1 >>
rect -4940 1810 -1820 1840
rect -4940 600 -3480 1810
rect -3430 600 -3370 1810
rect -3320 600 -3260 1810
rect -3210 600 -1820 1810
rect -4940 590 -1820 600
rect -4940 -880 -1820 -860
rect -4940 -2250 -4530 -880
rect -4480 -2250 -2910 -880
rect -2860 -2250 -2800 -880
rect -2750 -2250 -2690 -880
rect -2640 -2250 -1820 -880
rect -4940 -2260 -1820 -2250
rect -2150 -3370 -1820 -2260
rect -4930 -3400 -1820 -3370
rect -4930 -3450 -4700 -3400
rect -2360 -3450 -1820 -3400
rect -4930 -3510 -1820 -3450
rect -4930 -3560 -4700 -3510
rect -2360 -3560 -1820 -3510
rect -4930 -3620 -1820 -3560
rect -4930 -3670 -4700 -3620
rect -2360 -3670 -1820 -3620
rect -4930 -3700 -1820 -3670
rect -4930 -4350 -1820 -4320
rect -4930 -4400 -4700 -4350
rect -2360 -4400 -1820 -4350
rect -4930 -4460 -1820 -4400
rect -4930 -4510 -4700 -4460
rect -2360 -4510 -1820 -4460
rect -4930 -4570 -1820 -4510
rect -4930 -4620 -4700 -4570
rect -2360 -4620 -1820 -4570
rect -4930 -4990 -1820 -4620
rect -4930 -5040 -4700 -4990
rect -2360 -5040 -1820 -4990
rect -4930 -5170 -1820 -5040
rect -2020 -6070 -1820 -5170
rect -4940 -6080 -1820 -6070
rect -4940 -7460 -4540 -6080
rect -4490 -7460 -2920 -6080
rect -2870 -7460 -2810 -6080
rect -2760 -7460 -2700 -6080
rect -2650 -7460 -1820 -6080
rect -4940 -7470 -1820 -7460
rect -4940 -8950 -1820 -8940
rect -4940 -10180 -3490 -8950
rect -3440 -10180 -3380 -8950
rect -3330 -10180 -3270 -8950
rect -3220 -10180 -1820 -8950
rect -4940 -10190 -1820 -10180
<< labels >>
rlabel metal1 -4940 -9620 -4940 -9620 7 GND
rlabel metal1 -4940 -6810 -4940 -6810 7 VDD
rlabel metal1 -4940 -1560 -4940 -1560 7 GND
rlabel metal1 -4940 1060 -4940 1060 7 VDD
rlabel locali -4940 2480 -4940 2480 7 VCP
rlabel locali -4940 -11010 -4940 -11010 7 VCN
flabel locali -4930 -3200 -4930 -3200 0 FreeSans 640 0 0 0 VBN
port 1 nsew
rlabel locali -4940 -5410 -4940 -5410 7 VBP
port 2 w
<< end >>

magic
tech sky130A
timestamp 1702655834
<< locali >>
rect -60 1235 900 1255
rect -60 780 -40 1235
rect -20 1195 860 1215
rect -20 1030 0 1195
rect 840 1030 860 1195
rect 880 780 900 1235
rect -60 760 0 780
rect 840 760 900 780
use DFF  DFF_0
timestamp 1702606600
transform 1 0 -275 0 1 -295
box 695 295 1115 1500
use DFF  DFF_1
timestamp 1702606600
transform 1 0 -695 0 1 -295
box 695 295 1115 1500
<< end >>

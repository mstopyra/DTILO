magic
tech sky130A
timestamp 1702604723
<< nwell >>
rect -250 715 455 1775
<< nmos >>
rect -120 35 -105 635
rect 25 -365 40 635
rect 90 -365 105 635
rect 155 -365 170 635
rect 220 -365 235 635
rect 310 -15 325 635
<< pmos >>
rect -170 745 -155 1745
rect -105 745 -90 1745
rect 40 740 55 1740
rect 235 740 250 1740
rect 300 740 315 1740
rect 365 740 380 1740
<< ndiff >>
rect -170 620 -120 635
rect -170 50 -155 620
rect -135 50 -120 620
rect -170 35 -120 50
rect -105 620 -55 635
rect -105 50 -90 620
rect -70 50 -55 620
rect -105 35 -55 50
rect -25 620 25 635
rect -25 -350 -10 620
rect 10 -350 25 620
rect -25 -365 25 -350
rect 40 620 90 635
rect 40 -350 55 620
rect 75 -350 90 620
rect 40 -365 90 -350
rect 105 620 155 635
rect 105 -350 120 620
rect 140 -350 155 620
rect 105 -365 155 -350
rect 170 620 220 635
rect 170 -350 185 620
rect 205 -350 220 620
rect 170 -365 220 -350
rect 235 620 310 635
rect 235 -350 250 620
rect 270 -15 310 620
rect 325 620 375 635
rect 325 0 340 620
rect 360 0 375 620
rect 325 -15 375 0
rect 270 -350 285 -15
rect 235 -365 285 -350
<< pdiff >>
rect -220 1730 -170 1745
rect -220 760 -205 1730
rect -185 760 -170 1730
rect -220 745 -170 760
rect -155 1730 -105 1745
rect -155 760 -140 1730
rect -120 760 -105 1730
rect -155 745 -105 760
rect -90 1730 -40 1745
rect -90 760 -75 1730
rect -55 760 -40 1730
rect -90 745 -40 760
rect -10 1725 40 1740
rect -10 755 5 1725
rect 25 755 40 1725
rect -10 740 40 755
rect 55 1725 105 1740
rect 55 755 70 1725
rect 90 755 105 1725
rect 55 740 105 755
rect 190 1725 235 1740
rect 190 755 200 1725
rect 220 755 235 1725
rect 190 740 235 755
rect 250 1725 300 1740
rect 250 755 265 1725
rect 285 755 300 1725
rect 250 740 300 755
rect 315 1725 365 1740
rect 315 755 330 1725
rect 350 755 365 1725
rect 315 740 365 755
rect 380 1725 430 1740
rect 380 755 395 1725
rect 415 755 430 1725
rect 380 740 430 755
<< ndiffc >>
rect -155 50 -135 620
rect -90 50 -70 620
rect -10 -350 10 620
rect 55 -350 75 620
rect 120 -350 140 620
rect 185 -350 205 620
rect 250 -350 270 620
rect 340 0 360 620
<< pdiffc >>
rect -205 760 -185 1730
rect -140 760 -120 1730
rect -75 760 -55 1730
rect 5 755 25 1725
rect 70 755 90 1725
rect 200 755 220 1725
rect 265 755 285 1725
rect 330 755 350 1725
rect 395 755 415 1725
<< psubdiff >>
rect -220 620 -170 635
rect -220 50 -205 620
rect -185 50 -170 620
rect -220 35 -170 50
<< nsubdiff >>
rect 140 1725 190 1740
rect 140 755 155 1725
rect 175 755 190 1725
rect 140 740 190 755
<< psubdiffcont >>
rect -205 50 -185 620
<< nsubdiffcont >>
rect 155 755 175 1725
<< poly >>
rect 80 1785 120 1795
rect 80 1765 90 1785
rect 110 1770 120 1785
rect 110 1765 250 1770
rect -170 1745 -155 1760
rect -105 1745 -90 1760
rect 80 1755 250 1765
rect 40 1740 55 1755
rect 235 1740 250 1755
rect 300 1740 315 1755
rect 365 1740 380 1755
rect -170 730 -155 745
rect -105 730 -90 745
rect -255 710 -205 720
rect -255 680 -245 710
rect -215 705 -205 710
rect -170 715 -90 730
rect -55 715 -5 725
rect -170 705 -155 715
rect -215 685 -155 705
rect -215 680 -205 685
rect -255 670 -205 680
rect -120 635 -105 715
rect -55 685 -45 715
rect -15 705 -5 715
rect 40 705 55 740
rect 235 725 250 740
rect 300 725 315 740
rect 365 725 380 740
rect 235 710 380 725
rect -15 690 55 705
rect -15 685 -5 690
rect -55 675 -5 685
rect 40 665 55 690
rect 260 685 275 710
rect 260 670 325 685
rect 25 650 235 665
rect 25 635 40 650
rect 90 635 105 650
rect 155 635 170 650
rect 220 635 235 650
rect 310 635 325 670
rect -120 20 -105 35
rect 310 -30 325 -15
rect 25 -380 40 -365
rect 90 -380 105 -365
rect 155 -380 170 -365
rect 220 -380 235 -365
<< polycont >>
rect 90 1765 110 1785
rect -245 680 -215 710
rect -45 685 -15 715
<< locali >>
rect 80 1785 120 1795
rect -260 1760 -55 1780
rect -195 1740 -175 1760
rect -75 1740 -55 1760
rect 80 1765 90 1785
rect 110 1765 120 1785
rect 80 1755 120 1765
rect 210 1755 340 1775
rect -215 1730 -175 1740
rect -215 760 -205 1730
rect -185 760 -175 1730
rect -215 750 -175 760
rect -150 1730 -110 1740
rect -150 760 -140 1730
rect -120 760 -110 1730
rect -150 750 -110 760
rect -85 1730 -45 1740
rect 80 1735 100 1755
rect 210 1735 230 1755
rect 320 1735 340 1755
rect -85 760 -75 1730
rect -55 760 -45 1730
rect -85 750 -45 760
rect -5 1725 35 1735
rect -5 755 5 1725
rect 25 755 35 1725
rect -270 710 -205 720
rect -270 680 -245 710
rect -215 680 -205 710
rect -270 670 -205 680
rect -150 680 -130 750
rect -5 745 35 755
rect 60 1725 100 1735
rect 60 755 70 1725
rect 90 755 100 1725
rect 60 745 100 755
rect 145 1725 230 1735
rect 145 755 155 1725
rect 175 755 200 1725
rect 220 755 230 1725
rect 145 745 230 755
rect 255 1725 295 1735
rect 255 755 265 1725
rect 285 755 295 1725
rect 255 745 295 755
rect 320 1725 360 1735
rect 320 755 330 1725
rect 350 755 360 1725
rect 320 745 360 755
rect 385 1725 425 1735
rect 385 755 395 1725
rect 415 755 425 1725
rect 385 745 425 755
rect -55 715 -5 725
rect -55 700 -45 715
rect -100 685 -45 700
rect -15 685 -5 715
rect -100 680 -5 685
rect -150 660 -80 680
rect -55 675 -5 680
rect -100 630 -80 660
rect 60 670 80 745
rect 255 725 275 745
rect 385 725 405 745
rect 255 705 455 725
rect 60 650 195 670
rect 60 630 85 650
rect -215 620 -125 630
rect -215 50 -205 620
rect -185 50 -155 620
rect -135 50 -125 620
rect -215 40 -125 50
rect -100 620 -60 630
rect -100 50 -90 620
rect -70 50 -60 620
rect -100 0 -60 50
rect -20 620 20 630
rect -155 -100 -55 0
rect -20 -350 -10 620
rect 10 -350 20 620
rect -20 -360 20 -350
rect 45 620 85 630
rect 45 -350 55 620
rect 75 -350 85 620
rect 45 -360 85 -350
rect 110 620 150 630
rect 110 -350 120 620
rect 140 -350 150 620
rect 110 -360 150 -350
rect 175 625 195 650
rect 350 630 370 705
rect 430 660 455 705
rect 175 620 215 625
rect 175 -350 185 620
rect 205 -350 215 620
rect 175 -360 215 -350
rect 240 620 280 630
rect 240 -350 250 620
rect 270 -350 280 620
rect 330 620 370 630
rect 330 0 340 620
rect 360 0 370 620
rect 330 -10 370 0
rect 240 -360 280 -350
rect 0 -380 20 -360
rect 120 -380 140 -360
rect 240 -380 260 -360
rect 0 -400 260 -380
<< viali >>
rect 5 1100 25 1345
rect 200 1100 220 1345
rect -205 230 -185 470
rect -155 230 -135 470
rect -10 230 10 470
rect 250 230 270 470
<< metal1 >>
rect -255 1345 430 1350
rect -255 1100 5 1345
rect 25 1100 200 1345
rect 220 1100 430 1345
rect -255 1095 430 1100
rect -255 475 -220 480
rect -255 470 375 475
rect -255 230 -205 470
rect -185 230 -155 470
rect -135 230 -10 470
rect 10 230 250 470
rect 270 230 375 470
rect -255 225 375 230
rect -255 0 -240 225
rect -255 -15 -55 0
rect -155 -100 -55 -15
<< labels >>
flabel locali 455 715 455 715 0 FreeSans 400 0 0 0 Q
port 1 nsew
flabel locali -270 695 -270 695 0 FreeSans 400 0 0 0 A
port 2 nsew
flabel locali -260 1770 -260 1770 0 FreeSans 400 0 0 0 VP
port 3 nsew
flabel metal1 -255 1225 -255 1225 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 -155 -100 -55 0 0 FreeSans 360 0 0 0 C_L
flabel metal1 -255 340 -255 340 0 FreeSans 400 0 0 0 GND
port 5 nsew
<< end >>

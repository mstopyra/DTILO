magic
tech sky130A
timestamp 1702665350
<< nwell >>
rect -700 7700 17400 11100
<< nmos >>
rect 4800 3900 5200 7100
rect 5500 3900 5900 7100
rect 6800 3900 7200 7100
rect 7500 3900 7900 7100
rect 8800 3900 9200 7100
rect 9500 3900 9900 7100
rect 10800 3900 11200 7100
rect 11500 3900 11900 7100
rect 100 0 500 3200
rect 800 0 1200 3200
rect 2100 0 2500 3200
rect 2800 0 3200 3200
rect 4100 0 4500 3200
rect 4800 0 5200 3200
rect 6100 0 6500 3200
rect 6800 0 7200 3200
rect 7500 0 7900 3200
rect 8800 0 9200 3200
rect 9500 0 9900 3200
rect 10200 0 10600 3200
rect 11500 0 11900 3200
rect 12200 0 12600 3200
rect 13500 0 13900 3200
rect 14200 0 14600 3200
rect 15500 0 15900 3200
rect 16200 0 16600 3200
<< pmos >>
rect 3500 7800 3900 11000
rect 4200 7800 4600 11000
rect 5500 7800 5900 11000
rect 6200 7800 6600 11000
rect 7500 7800 7900 11000
rect 8800 7800 9200 11000
rect 10100 7800 10500 11000
rect 10800 7800 11200 11000
rect 12100 7800 12500 11000
rect 12800 7800 13200 11000
<< ndiff >>
rect 4500 7000 4800 7100
rect 4500 4000 4600 7000
rect 4700 4000 4800 7000
rect 4500 3900 4800 4000
rect 5200 7000 5500 7100
rect 5200 4000 5300 7000
rect 5400 4000 5500 7000
rect 5200 3900 5500 4000
rect 5900 7000 6200 7100
rect 6500 7000 6800 7100
rect 5900 4000 6000 7000
rect 6100 4000 6200 7000
rect 6500 4000 6600 7000
rect 6700 4000 6800 7000
rect 5900 3900 6200 4000
rect 6500 3900 6800 4000
rect 7200 7000 7500 7100
rect 7200 4000 7300 7000
rect 7400 4000 7500 7000
rect 7200 3900 7500 4000
rect 7900 7000 8200 7100
rect 8500 7000 8800 7100
rect 7900 4000 8000 7000
rect 8100 4000 8200 7000
rect 8500 4000 8600 7000
rect 8700 4000 8800 7000
rect 7900 3900 8200 4000
rect 8500 3900 8800 4000
rect 9200 7000 9500 7100
rect 9200 4000 9300 7000
rect 9400 4000 9500 7000
rect 9200 3900 9500 4000
rect 9900 7000 10200 7100
rect 10500 7000 10800 7100
rect 9900 4000 10000 7000
rect 10100 4000 10200 7000
rect 10500 4000 10600 7000
rect 10700 4000 10800 7000
rect 9900 3900 10200 4000
rect 10500 3900 10800 4000
rect 11200 7000 11500 7100
rect 11200 4000 11300 7000
rect 11400 4000 11500 7000
rect 11200 3900 11500 4000
rect 11900 7000 12200 7100
rect 11900 4000 12000 7000
rect 12100 4000 12200 7000
rect 11900 3900 12200 4000
rect -200 3100 100 3200
rect -200 100 -100 3100
rect 0 100 100 3100
rect -200 0 100 100
rect 500 3100 800 3200
rect 500 100 600 3100
rect 700 100 800 3100
rect 500 0 800 100
rect 1200 3100 1500 3200
rect 1800 3100 2100 3200
rect 1200 100 1300 3100
rect 1400 100 1500 3100
rect 1800 100 1900 3100
rect 2000 100 2100 3100
rect 1200 0 1500 100
rect 1800 0 2100 100
rect 2500 3100 2800 3200
rect 2500 100 2600 3100
rect 2700 100 2800 3100
rect 2500 0 2800 100
rect 3200 3100 3500 3200
rect 3800 3100 4100 3200
rect 3200 100 3300 3100
rect 3400 100 3500 3100
rect 3800 100 3900 3100
rect 4000 100 4100 3100
rect 3200 0 3500 100
rect 3800 0 4100 100
rect 4500 3100 4800 3200
rect 4500 100 4600 3100
rect 4700 100 4800 3100
rect 4500 0 4800 100
rect 5200 3100 5500 3200
rect 5800 3100 6100 3200
rect 5200 100 5300 3100
rect 5400 100 5500 3100
rect 5800 100 5900 3100
rect 6000 100 6100 3100
rect 5200 0 5500 100
rect 5800 0 6100 100
rect 6500 3100 6800 3200
rect 6500 100 6600 3100
rect 6700 100 6800 3100
rect 6500 0 6800 100
rect 7200 3100 7500 3200
rect 7200 100 7300 3100
rect 7400 100 7500 3100
rect 7200 0 7500 100
rect 7900 3100 8200 3200
rect 8500 3100 8800 3200
rect 7900 100 8000 3100
rect 8100 100 8200 3100
rect 8500 100 8600 3100
rect 8700 100 8800 3100
rect 7900 0 8200 100
rect 8500 0 8800 100
rect 9200 3100 9500 3200
rect 9200 100 9300 3100
rect 9400 100 9500 3100
rect 9200 0 9500 100
rect 9900 3100 10200 3200
rect 9900 100 10000 3100
rect 10100 100 10200 3100
rect 9900 0 10200 100
rect 10600 3100 10900 3200
rect 11200 3100 11500 3200
rect 10600 100 10700 3100
rect 10800 100 10900 3100
rect 11200 100 11300 3100
rect 11400 100 11500 3100
rect 10600 0 10900 100
rect 11200 0 11500 100
rect 11900 3100 12200 3200
rect 11900 100 12000 3100
rect 12100 100 12200 3100
rect 11900 0 12200 100
rect 12600 3100 12900 3200
rect 13200 3100 13500 3200
rect 12600 100 12700 3100
rect 12800 100 12900 3100
rect 13200 100 13300 3100
rect 13400 100 13500 3100
rect 12600 0 12900 100
rect 13200 0 13500 100
rect 13900 3100 14200 3200
rect 13900 100 14000 3100
rect 14100 100 14200 3100
rect 13900 0 14200 100
rect 14600 3100 14900 3200
rect 15200 3100 15500 3200
rect 14600 100 14700 3100
rect 14800 100 14900 3100
rect 15200 100 15300 3100
rect 15400 100 15500 3100
rect 14600 0 14900 100
rect 15200 0 15500 100
rect 15900 3100 16200 3200
rect 15900 100 16000 3100
rect 16100 100 16200 3100
rect 15900 0 16200 100
rect 16600 3100 16900 3200
rect 16600 100 16700 3100
rect 16800 100 16900 3100
rect 16600 0 16900 100
<< pdiff >>
rect 3200 10900 3500 11000
rect 3200 7900 3300 10900
rect 3400 7900 3500 10900
rect 3200 7800 3500 7900
rect 3900 10900 4200 11000
rect 3900 7900 4000 10900
rect 4100 7900 4200 10900
rect 3900 7800 4200 7900
rect 4600 10900 4900 11000
rect 5200 10900 5500 11000
rect 4600 7900 4700 10900
rect 4800 7900 4900 10900
rect 5200 7900 5300 10900
rect 5400 7900 5500 10900
rect 4600 7800 4900 7900
rect 5200 7800 5500 7900
rect 5900 10900 6200 11000
rect 5900 7900 6000 10900
rect 6100 7900 6200 10900
rect 5900 7800 6200 7900
rect 6600 10900 6900 11000
rect 7200 10900 7500 11000
rect 6600 7900 6700 10900
rect 6800 7900 6900 10900
rect 7200 7900 7300 10900
rect 7400 7900 7500 10900
rect 6600 7800 6900 7900
rect 7200 7800 7500 7900
rect 7900 10900 8200 11000
rect 8500 10900 8800 11000
rect 7900 7900 8000 10900
rect 8100 7900 8200 10900
rect 8500 7900 8600 10900
rect 8700 7900 8800 10900
rect 7900 7800 8200 7900
rect 8500 7800 8800 7900
rect 9200 10900 9500 11000
rect 9800 10900 10100 11000
rect 9200 7900 9300 10900
rect 9400 7900 9500 10900
rect 9800 7900 9900 10900
rect 10000 7900 10100 10900
rect 9200 7800 9500 7900
rect 9800 7800 10100 7900
rect 10500 10900 10800 11000
rect 10500 7900 10600 10900
rect 10700 7900 10800 10900
rect 10500 7800 10800 7900
rect 11200 10900 11500 11000
rect 11800 10900 12100 11000
rect 11200 7900 11300 10900
rect 11400 7900 11500 10900
rect 11800 7900 11900 10900
rect 12000 7900 12100 10900
rect 11200 7800 11500 7900
rect 11800 7800 12100 7900
rect 12500 10900 12800 11000
rect 12500 7900 12600 10900
rect 12700 7900 12800 10900
rect 12500 7800 12800 7900
rect 13200 10900 13500 11000
rect 13200 7900 13300 10900
rect 13400 7900 13500 10900
rect 13200 7800 13500 7900
<< ndiffc >>
rect 4600 4000 4700 7000
rect 5300 4000 5400 7000
rect 6000 4000 6100 7000
rect 6600 4000 6700 7000
rect 7300 4000 7400 7000
rect 8000 4000 8100 7000
rect 8600 4000 8700 7000
rect 9300 4000 9400 7000
rect 10000 4000 10100 7000
rect 10600 4000 10700 7000
rect 11300 4000 11400 7000
rect 12000 4000 12100 7000
rect -100 100 0 3100
rect 600 100 700 3100
rect 1300 100 1400 3100
rect 1900 100 2000 3100
rect 2600 100 2700 3100
rect 3300 100 3400 3100
rect 3900 100 4000 3100
rect 4600 100 4700 3100
rect 5300 100 5400 3100
rect 5900 100 6000 3100
rect 6600 100 6700 3100
rect 7300 100 7400 3100
rect 8000 100 8100 3100
rect 8600 100 8700 3100
rect 9300 100 9400 3100
rect 10000 100 10100 3100
rect 10700 100 10800 3100
rect 11300 100 11400 3100
rect 12000 100 12100 3100
rect 12700 100 12800 3100
rect 13300 100 13400 3100
rect 14000 100 14100 3100
rect 14700 100 14800 3100
rect 15300 100 15400 3100
rect 16000 100 16100 3100
rect 16700 100 16800 3100
<< pdiffc >>
rect 3300 7900 3400 10900
rect 4000 7900 4100 10900
rect 4700 7900 4800 10900
rect 5300 7900 5400 10900
rect 6000 7900 6100 10900
rect 6700 7900 6800 10900
rect 7300 7900 7400 10900
rect 8000 7900 8100 10900
rect 8600 7900 8700 10900
rect 9300 7900 9400 10900
rect 9900 7900 10000 10900
rect 10600 7900 10700 10900
rect 11300 7900 11400 10900
rect 11900 7900 12000 10900
rect 12600 7900 12700 10900
rect 13300 7900 13400 10900
<< psubdiff >>
rect 4200 7000 4500 7100
rect 4200 4000 4300 7000
rect 4400 4000 4500 7000
rect 4200 3900 4500 4000
rect 6200 7000 6500 7100
rect 6200 4000 6300 7000
rect 6400 4000 6500 7000
rect 6200 3900 6500 4000
rect 8200 7000 8500 7100
rect 8200 4000 8300 7000
rect 8400 4000 8500 7000
rect 8200 3900 8500 4000
rect 10200 7000 10500 7100
rect 10200 4000 10300 7000
rect 10400 4000 10500 7000
rect 10200 3900 10500 4000
rect 12200 7000 12500 7100
rect 12200 4000 12300 7000
rect 12400 4000 12500 7000
rect 12200 3900 12500 4000
rect -500 3100 -200 3200
rect -500 100 -400 3100
rect -300 100 -200 3100
rect -500 0 -200 100
rect 1500 3100 1800 3200
rect 1500 100 1600 3100
rect 1700 100 1800 3100
rect 1500 0 1800 100
rect 3500 3100 3800 3200
rect 3500 100 3600 3100
rect 3700 100 3800 3100
rect 3500 0 3800 100
rect 5500 3100 5800 3200
rect 5500 100 5600 3100
rect 5700 100 5800 3100
rect 5500 0 5800 100
rect 8200 3100 8500 3200
rect 8200 100 8300 3100
rect 8400 100 8500 3100
rect 8200 0 8500 100
rect 10900 3100 11200 3200
rect 10900 100 11000 3100
rect 11100 100 11200 3100
rect 10900 0 11200 100
rect 12900 3100 13200 3200
rect 12900 100 13000 3100
rect 13100 100 13200 3100
rect 12900 0 13200 100
rect 14900 3100 15200 3200
rect 14900 100 15000 3100
rect 15100 100 15200 3100
rect 14900 0 15200 100
rect 16900 3100 17200 3200
rect 16900 100 17000 3100
rect 17100 100 17200 3100
rect 16900 0 17200 100
<< nsubdiff >>
rect 2900 10900 3200 11000
rect 2900 7900 3000 10900
rect 3100 7900 3200 10900
rect 2900 7800 3200 7900
rect 4900 10900 5200 11000
rect 4900 7900 5000 10900
rect 5100 7900 5200 10900
rect 4900 7800 5200 7900
rect 6900 10900 7200 11000
rect 6900 7900 7000 10900
rect 7100 7900 7200 10900
rect 6900 7800 7200 7900
rect 8200 10900 8500 11000
rect 8200 7900 8300 10900
rect 8400 7900 8500 10900
rect 8200 7800 8500 7900
rect 9500 10900 9800 11000
rect 9500 7900 9600 10900
rect 9700 7900 9800 10900
rect 9500 7800 9800 7900
rect 11500 10900 11800 11000
rect 11500 7900 11600 10900
rect 11700 7900 11800 10900
rect 11500 7800 11800 7900
rect 13500 10900 13800 11000
rect 13500 7900 13600 10900
rect 13700 7900 13800 10900
rect 13500 7800 13800 7900
<< psubdiffcont >>
rect 4300 4000 4400 7000
rect 6300 4000 6400 7000
rect 8300 4000 8400 7000
rect 10300 4000 10400 7000
rect 12300 4000 12400 7000
rect -400 100 -300 3100
rect 1600 100 1700 3100
rect 3600 100 3700 3100
rect 5600 100 5700 3100
rect 8300 100 8400 3100
rect 11000 100 11100 3100
rect 13000 100 13100 3100
rect 15000 100 15100 3100
rect 17000 100 17100 3100
<< nsubdiffcont >>
rect 3000 7900 3100 10900
rect 5000 7900 5100 10900
rect 7000 7900 7100 10900
rect 8300 7900 8400 10900
rect 9600 7900 9700 10900
rect 11600 7900 11700 10900
rect 13600 7900 13700 10900
<< poly >>
rect 3500 11000 3900 11100
rect 4200 11000 4600 11100
rect 5500 11000 5900 11100
rect 6200 11000 6600 11100
rect 7500 11000 7900 11100
rect 8800 11000 9200 11100
rect 10100 11000 10500 11100
rect 10800 11000 11200 11100
rect 12100 11000 12500 11100
rect 12800 11000 13200 11100
rect 3500 7650 3900 7800
rect 3500 7550 3550 7650
rect 3850 7550 3900 7650
rect 3500 7500 3900 7550
rect 4200 7500 4600 7800
rect 5500 7750 5900 7800
rect 5500 7650 5550 7750
rect 5850 7700 5900 7750
rect 6200 7700 6600 7800
rect 5850 7650 6600 7700
rect 5500 7600 6600 7650
rect 7500 7650 7900 7800
rect 6700 7550 6900 7600
rect 6700 7500 6750 7550
rect 4200 7450 6750 7500
rect 6850 7500 6900 7550
rect 7500 7500 7550 7650
rect 6850 7450 7550 7500
rect 7850 7500 7900 7650
rect 8800 7500 9200 7800
rect 10100 7700 10500 7800
rect 10800 7750 11200 7800
rect 10800 7700 10850 7750
rect 10100 7650 10850 7700
rect 11150 7650 11200 7750
rect 10100 7600 11200 7650
rect 9800 7550 10000 7600
rect 9800 7500 9850 7550
rect 7850 7450 9850 7500
rect 9950 7500 10000 7550
rect 12100 7500 12500 7800
rect 12800 7650 13200 7800
rect 12800 7550 12850 7650
rect 13150 7550 13200 7650
rect 12800 7500 13200 7550
rect 9950 7450 12500 7500
rect 4200 7400 12500 7450
rect 4800 7100 5200 7200
rect 5500 7100 5900 7200
rect 6800 7100 7200 7200
rect 7500 7100 7900 7200
rect 8800 7100 9200 7200
rect 9500 7100 9900 7200
rect 10800 7100 11200 7200
rect 11500 7100 11900 7200
rect 4800 3850 5200 3900
rect 4800 3750 4850 3850
rect 5150 3750 5200 3850
rect 5500 3800 5900 3900
rect 4800 3700 5200 3750
rect 5800 3400 5900 3800
rect 6800 3800 7200 3900
rect 7500 3850 7900 3900
rect 7500 3800 7550 3850
rect 6800 3750 7550 3800
rect 7850 3750 7900 3850
rect 6800 3700 7900 3750
rect 8800 3850 9200 3900
rect 8800 3650 8850 3850
rect 9150 3800 9200 3850
rect 9500 3800 9900 3900
rect 9150 3700 9900 3800
rect 10800 3800 11200 3900
rect 11500 3850 11900 3900
rect 9150 3650 9200 3700
rect 8800 3600 9200 3650
rect 10800 3400 10900 3800
rect 11500 3750 11550 3850
rect 11850 3750 11900 3850
rect 11500 3700 11900 3750
rect 5800 3300 6200 3400
rect 10500 3300 10900 3400
rect 100 3200 500 3300
rect 800 3200 1200 3300
rect 2100 3200 2500 3300
rect 2800 3200 3200 3300
rect 4100 3200 4500 3300
rect 4800 3200 5200 3300
rect 6100 3200 6500 3300
rect 6800 3200 7200 3300
rect 7500 3200 7900 3300
rect 8800 3200 9200 3300
rect 9500 3200 9900 3300
rect 10200 3200 10600 3300
rect 11500 3200 11900 3300
rect 12200 3200 12600 3300
rect 13500 3200 13900 3300
rect 14200 3200 14600 3300
rect 15500 3200 15900 3300
rect 16200 3200 16600 3300
rect 100 -150 500 0
rect 800 -100 1200 0
rect 2100 -100 2500 0
rect 2800 -100 3200 0
rect 4100 -100 4500 0
rect 4800 -100 5200 0
rect 6100 -100 6500 0
rect 6800 -100 7200 0
rect 7500 -100 7900 0
rect 8800 -100 9200 0
rect 9500 -100 9900 0
rect 10200 -100 10600 0
rect 11500 -100 11900 0
rect 12200 -100 12600 0
rect 13500 -100 13900 0
rect 14200 -100 14600 0
rect 15500 -100 15900 0
rect 100 -250 150 -150
rect 450 -250 500 -150
rect 100 -300 500 -250
rect 600 -150 8100 -100
rect 600 -250 650 -150
rect 750 -250 1250 -150
rect 1450 -250 1850 -150
rect 2050 -250 2550 -150
rect 2750 -250 3250 -150
rect 3450 -250 3850 -150
rect 4050 -250 4550 -150
rect 4750 -250 5250 -150
rect 5450 -250 5850 -150
rect 6050 -250 6550 -150
rect 6750 -250 7250 -150
rect 7450 -250 7950 -150
rect 8050 -250 8100 -150
rect 600 -300 8100 -250
rect 8600 -150 16100 -100
rect 8600 -250 8650 -150
rect 8750 -250 9250 -150
rect 9450 -250 9950 -150
rect 10150 -250 10650 -150
rect 10850 -250 11250 -150
rect 11450 -250 11950 -150
rect 12150 -250 12650 -150
rect 12850 -250 13250 -150
rect 13450 -250 13950 -150
rect 14150 -250 14650 -150
rect 14850 -250 15250 -150
rect 15450 -250 15950 -150
rect 16050 -250 16100 -150
rect 8600 -300 16100 -250
rect 16200 -150 16600 0
rect 16200 -250 16250 -150
rect 16550 -250 16600 -150
rect 16200 -300 16600 -250
<< polycont >>
rect 3550 7550 3850 7650
rect 5550 7650 5850 7750
rect 6750 7450 6850 7550
rect 7550 7450 7850 7650
rect 10850 7650 11150 7750
rect 9850 7450 9950 7550
rect 12850 7550 13150 7650
rect 4850 3750 5150 3850
rect 7550 3750 7850 3850
rect 8850 3650 9150 3850
rect 11550 3750 11850 3850
rect 150 -250 450 -150
rect 650 -250 750 -150
rect 1250 -250 1450 -150
rect 1850 -250 2050 -150
rect 2550 -250 2750 -150
rect 3250 -250 3450 -150
rect 3850 -250 4050 -150
rect 4550 -250 4750 -150
rect 5250 -250 5450 -150
rect 5850 -250 6050 -150
rect 6550 -250 6750 -150
rect 7250 -250 7450 -150
rect 7950 -250 8050 -150
rect 8650 -250 8750 -150
rect 9250 -250 9450 -150
rect 9950 -250 10150 -150
rect 10650 -250 10850 -150
rect 11250 -250 11450 -150
rect 11950 -250 12150 -150
rect 12650 -250 12850 -150
rect 13250 -250 13450 -150
rect 13950 -250 14150 -150
rect 14650 -250 14850 -150
rect 15250 -250 15450 -150
rect 15950 -250 16050 -150
rect 16250 -250 16550 -150
<< locali >>
rect 3000 10900 3100 11000
rect 3300 10900 3400 11000
rect 5000 10900 5100 11000
rect 6000 10900 6100 11000
rect 7000 10900 7100 11000
rect 7300 10900 7400 11000
rect 8300 10900 8400 11000
rect 9300 10900 9400 11000
rect 9600 10900 9700 11000
rect 10600 10900 10700 11000
rect 11600 10900 11700 11000
rect 13300 10900 13400 11000
rect 13600 10900 13700 11000
rect 3100 7900 3300 10900
rect 3400 7900 3500 10900
rect 3900 7900 4000 10900
rect 4100 7900 4200 10900
rect 4600 7900 4700 10900
rect 4800 7900 4900 10900
rect 5200 7900 5300 10900
rect 5400 7900 5500 10900
rect 5900 7900 6000 10900
rect 6100 7900 6200 10900
rect 6600 7900 6700 10900
rect 6800 7900 6900 10900
rect 7200 7900 7300 10900
rect 7400 7900 7500 10900
rect 7900 7900 8000 10900
rect 8100 7900 8200 10900
rect 8500 7900 8600 10900
rect 8700 7900 8800 10900
rect 9200 7900 9300 10900
rect 9400 7900 9500 10900
rect 9800 7900 9900 10900
rect 10000 7900 10100 10900
rect 10500 7900 10600 10900
rect 10700 7900 10800 10900
rect 11200 7900 11300 10900
rect 11400 7900 11500 10900
rect 11800 7900 11900 10900
rect 12000 7900 12100 10900
rect 12500 7900 12600 10900
rect 12700 7900 12800 10900
rect 13200 7900 13300 10900
rect 13400 7900 13600 10900
rect 3000 7800 3100 7900
rect 3300 7650 3400 7900
rect 3500 7650 3900 7700
rect 3300 7550 3550 7650
rect 3850 7550 3900 7650
rect 3500 7500 3900 7550
rect 4000 3850 4100 7900
rect 5000 7800 5100 7900
rect 5300 7700 5400 7900
rect 5500 7750 5900 7800
rect 5500 7700 5550 7750
rect 5300 7650 5550 7700
rect 5850 7650 5900 7750
rect 5300 7600 5900 7650
rect 6700 7600 6800 7900
rect 7000 7800 7100 7900
rect 7500 7650 7900 7700
rect 4300 7000 4400 7100
rect 5300 7000 5400 7600
rect 6700 7550 6900 7600
rect 6700 7500 6750 7550
rect 6600 7450 6750 7500
rect 6850 7450 6900 7550
rect 6600 7400 6900 7450
rect 7500 7450 7550 7650
rect 7850 7450 7900 7650
rect 7500 7400 7900 7450
rect 6300 7000 6400 7100
rect 6600 7000 6700 7400
rect 8000 7000 8100 7900
rect 8300 7800 8400 7900
rect 8300 7000 8400 7100
rect 8600 7000 8700 7900
rect 9600 7800 9700 7900
rect 9900 7600 10000 7900
rect 10800 7750 11200 7800
rect 10800 7650 10850 7750
rect 11150 7700 11200 7750
rect 11300 7700 11400 7900
rect 11600 7800 11700 7900
rect 11150 7650 11400 7700
rect 10800 7600 11400 7650
rect 9800 7550 10000 7600
rect 9800 7450 9850 7550
rect 9950 7500 10000 7550
rect 9950 7450 10100 7500
rect 9800 7400 10100 7450
rect 10000 7000 10100 7400
rect 10300 7000 10400 7100
rect 11300 7000 11400 7600
rect 12300 7000 12400 7100
rect 4400 4000 4600 7000
rect 4700 4000 4800 7000
rect 5200 4000 5300 7000
rect 5400 4000 5500 7000
rect 5900 4000 6000 7000
rect 6100 4000 6200 7000
rect 6500 4000 6600 7000
rect 6700 4000 6800 7000
rect 7200 4000 7300 7000
rect 7400 4000 7500 7000
rect 7900 4000 8000 7000
rect 8100 4000 8200 7000
rect 8500 4000 8600 7000
rect 8700 4000 8800 7000
rect 9200 4000 9300 7000
rect 9400 4000 9500 7000
rect 9900 4000 10000 7000
rect 10100 4000 10200 7000
rect 10500 4000 10600 7000
rect 10700 4000 10800 7000
rect 11200 4000 11300 7000
rect 11400 4000 11500 7000
rect 11900 4000 12000 7000
rect 12100 4000 12300 7000
rect 4300 3900 4400 4000
rect -100 3750 4100 3850
rect 4600 3850 4700 4000
rect 4800 3850 5200 3900
rect 4600 3750 4850 3850
rect 5150 3750 5200 3850
rect -400 3100 -300 3200
rect -100 3100 0 3750
rect 4800 3700 5200 3750
rect 6000 3700 6100 4000
rect 6300 3900 6400 4000
rect 7300 3700 7400 4000
rect 7500 3850 7900 3900
rect 7500 3750 7550 3850
rect 7850 3800 7900 3850
rect 8000 3800 8100 4000
rect 8300 3900 8400 4000
rect 8600 3800 8700 4000
rect 8800 3850 9200 3900
rect 8800 3800 8850 3850
rect 7850 3750 8850 3800
rect 7500 3700 8850 3750
rect 6000 3650 7400 3700
rect 6000 3600 6250 3650
rect 6200 3450 6250 3600
rect 6450 3600 7400 3650
rect 8800 3650 8850 3700
rect 9150 3650 9200 3850
rect 8800 3600 9200 3650
rect 9300 3700 9400 4000
rect 10300 3900 10400 4000
rect 10600 3700 10700 4000
rect 11500 3850 11900 3900
rect 12000 3850 12100 4000
rect 12300 3900 12400 4000
rect 11500 3750 11550 3850
rect 11850 3750 12100 3850
rect 12600 3850 12700 7900
rect 12800 7650 13200 7700
rect 13300 7650 13400 7900
rect 13600 7800 13700 7900
rect 12800 7550 12850 7650
rect 13150 7550 13400 7650
rect 12800 7500 13200 7550
rect 12600 3750 16800 3850
rect 11500 3700 11900 3750
rect 9300 3650 10700 3700
rect 9300 3600 10250 3650
rect 6450 3450 6500 3600
rect 6200 3400 6500 3450
rect 10200 3450 10250 3600
rect 10450 3600 10700 3650
rect 10450 3450 10500 3600
rect 10200 3400 10500 3450
rect 1600 3100 1700 3200
rect 3600 3100 3700 3200
rect 5600 3100 5700 3200
rect 8300 3100 8400 3200
rect 11000 3100 11100 3200
rect 13000 3100 13100 3200
rect 15000 3100 15100 3200
rect 16700 3100 16800 3750
rect 17000 3100 17100 3200
rect -300 100 -100 3100
rect 0 100 100 3100
rect 500 100 600 3100
rect 700 100 800 3100
rect 1200 100 1300 3100
rect 1400 100 1500 3100
rect 1800 100 1900 3100
rect 2000 100 2100 3100
rect 2500 100 2600 3100
rect 2700 100 2800 3100
rect 3200 100 3300 3100
rect 3400 100 3500 3100
rect 3800 100 3900 3100
rect 4000 100 4100 3100
rect 4500 100 4600 3100
rect 4700 100 4800 3100
rect 5200 100 5300 3100
rect 5400 100 5500 3100
rect 5800 100 5900 3100
rect 6000 100 6100 3100
rect 6500 100 6600 3100
rect 6700 100 6800 3100
rect 7200 100 7300 3100
rect 7400 100 7500 3100
rect 7900 100 8000 3100
rect 8100 100 8200 3100
rect 8500 100 8600 3100
rect 8700 100 8800 3100
rect 9200 100 9300 3100
rect 9400 100 9500 3100
rect 9900 100 10000 3100
rect 10100 100 10200 3100
rect 10600 100 10700 3100
rect 10800 100 10900 3100
rect 11200 100 11300 3100
rect 11400 100 11500 3100
rect 11900 100 12000 3100
rect 12100 100 12200 3100
rect 12600 100 12700 3100
rect 12800 100 12900 3100
rect 13200 100 13300 3100
rect 13400 100 13500 3100
rect 13900 100 14000 3100
rect 14100 100 14200 3100
rect 14600 100 14700 3100
rect 14800 100 14900 3100
rect 15200 100 15300 3100
rect 15400 100 15500 3100
rect 15900 100 16000 3100
rect 16100 100 16200 3100
rect 16600 100 16700 3100
rect 16800 100 17000 3100
rect -400 0 100 100
rect -100 -150 0 0
rect 600 -100 700 100
rect 1300 -100 1400 100
rect 1600 0 1700 100
rect 1900 -100 2000 100
rect 2600 -100 2700 100
rect 3300 -100 3400 100
rect 3600 0 3700 100
rect 3900 -100 4000 100
rect 4600 -100 4700 100
rect 5300 -100 5400 100
rect 5600 0 5700 100
rect 5900 -100 6000 100
rect 6600 -100 6700 100
rect 7300 -100 7400 100
rect 8000 -100 8100 100
rect 8300 0 8400 100
rect 100 -150 500 -100
rect -100 -250 150 -150
rect 450 -250 500 -150
rect 100 -300 500 -250
rect 600 -150 800 -100
rect 600 -250 650 -150
rect 750 -250 800 -150
rect 600 -300 800 -250
rect 1200 -150 1500 -100
rect 1200 -250 1250 -150
rect 1450 -250 1500 -150
rect 1200 -300 1500 -250
rect 1800 -150 2100 -100
rect 1800 -250 1850 -150
rect 2050 -250 2100 -150
rect 1800 -300 2100 -250
rect 2500 -150 2800 -100
rect 2500 -250 2550 -150
rect 2750 -250 2800 -150
rect 2500 -300 2800 -250
rect 3200 -150 3500 -100
rect 3200 -250 3250 -150
rect 3450 -250 3500 -150
rect 3200 -300 3500 -250
rect 3800 -150 4100 -100
rect 3800 -250 3850 -150
rect 4050 -250 4100 -150
rect 3800 -300 4100 -250
rect 4500 -150 4800 -100
rect 4500 -250 4550 -150
rect 4750 -250 4800 -150
rect 4500 -300 4800 -250
rect 5200 -150 5500 -100
rect 5200 -250 5250 -150
rect 5450 -250 5500 -150
rect 5200 -300 5500 -250
rect 5800 -150 6100 -100
rect 5800 -250 5850 -150
rect 6050 -250 6100 -150
rect 5800 -300 6100 -250
rect 6500 -150 6800 -100
rect 6500 -250 6550 -150
rect 6750 -250 6800 -150
rect 6500 -300 6800 -250
rect 7200 -150 7500 -100
rect 7200 -250 7250 -150
rect 7450 -250 7500 -150
rect 7200 -300 7500 -250
rect 7900 -150 8100 -100
rect 7900 -250 7950 -150
rect 8050 -250 8100 -150
rect 7900 -300 8100 -250
rect 8600 -100 8700 100
rect 9300 -100 9400 100
rect 10000 -100 10100 100
rect 10700 -100 10800 100
rect 11000 0 11100 100
rect 11300 -100 11400 100
rect 12000 -100 12100 100
rect 12700 -100 12800 100
rect 13000 0 13100 100
rect 13300 -100 13400 100
rect 14000 -100 14100 100
rect 14700 -100 14800 100
rect 15000 0 15100 100
rect 15300 -100 15400 100
rect 16000 -100 16100 100
rect 16600 0 17100 100
rect 8600 -150 8800 -100
rect 8600 -250 8650 -150
rect 8750 -250 8800 -150
rect 8600 -300 8800 -250
rect 9200 -150 9500 -100
rect 9200 -250 9250 -150
rect 9450 -250 9500 -150
rect 9200 -300 9500 -250
rect 9900 -150 10200 -100
rect 9900 -250 9950 -150
rect 10150 -250 10200 -150
rect 9900 -300 10200 -250
rect 10600 -150 10900 -100
rect 10600 -250 10650 -150
rect 10850 -250 10900 -150
rect 10600 -300 10900 -250
rect 11200 -150 11500 -100
rect 11200 -250 11250 -150
rect 11450 -250 11500 -150
rect 11200 -300 11500 -250
rect 11900 -150 12200 -100
rect 11900 -250 11950 -150
rect 12150 -250 12200 -150
rect 11900 -300 12200 -250
rect 12600 -150 12900 -100
rect 12600 -250 12650 -150
rect 12850 -250 12900 -150
rect 12600 -300 12900 -250
rect 13200 -150 13500 -100
rect 13200 -250 13250 -150
rect 13450 -250 13500 -150
rect 13200 -300 13500 -250
rect 13900 -150 14200 -100
rect 13900 -250 13950 -150
rect 14150 -250 14200 -150
rect 13900 -300 14200 -250
rect 14600 -150 14900 -100
rect 14600 -250 14650 -150
rect 14850 -250 14900 -150
rect 14600 -300 14900 -250
rect 15200 -150 15500 -100
rect 15200 -250 15250 -150
rect 15450 -250 15500 -150
rect 15200 -300 15500 -250
rect 15900 -150 16100 -100
rect 15900 -250 15950 -150
rect 16050 -250 16100 -150
rect 15900 -300 16100 -250
rect 16200 -150 16600 -100
rect 16700 -150 16800 0
rect 16200 -250 16250 -150
rect 16550 -250 16800 -150
rect 16200 -300 16600 -250
<< viali >>
rect 3000 7900 3100 10900
rect 5000 7900 5100 10900
rect 6000 7900 6100 10900
rect 7000 7900 7100 10900
rect 7300 7900 7400 10900
rect 8300 7900 8400 10900
rect 9300 7900 9400 10900
rect 9600 7900 9700 10900
rect 10600 7900 10700 10900
rect 11600 7900 11700 10900
rect 13600 7900 13700 10900
rect 7550 7450 7850 7650
rect 4300 4000 4400 7000
rect 6300 4000 6400 7000
rect 8300 4000 8400 7000
rect 10300 4000 10400 7000
rect 12300 4000 12400 7000
rect 6250 3450 6450 3650
rect 8850 3650 9150 3850
rect 10250 3450 10450 3650
rect -400 100 -300 3100
rect 1600 100 1700 3100
rect 3600 100 3700 3100
rect 5600 100 5700 3100
rect 8300 100 8400 3100
rect 11000 100 11100 3100
rect 13000 100 13100 3100
rect 15000 100 15100 3100
rect 17000 100 17100 3100
<< metal1 >>
rect -700 10900 17400 11000
rect -700 7900 3000 10900
rect 3100 7900 5000 10900
rect 5100 7900 6000 10900
rect 6100 7900 7000 10900
rect 7100 7900 7300 10900
rect 7400 7900 8300 10900
rect 8400 7900 9300 10900
rect 9400 7900 9600 10900
rect 9700 7900 10600 10900
rect 10700 7900 11600 10900
rect 11700 7900 13600 10900
rect 13700 7900 17400 10900
rect -700 7800 17400 7900
rect 7500 7650 7900 7700
rect 7500 7450 7550 7650
rect 7850 7450 7900 7650
rect 7500 7400 7900 7450
rect 4200 7000 4500 7100
rect 4200 4000 4300 7000
rect 4400 4000 4500 7000
rect 4200 3200 4500 4000
rect 6200 7000 6500 7100
rect 6200 4000 6300 7000
rect 6400 4000 6500 7000
rect 6200 3650 6500 4000
rect 6200 3450 6250 3650
rect 6450 3450 6500 3650
rect 6200 3200 6500 3450
rect 8200 7000 8500 7100
rect 8200 4000 8300 7000
rect 8400 4000 8500 7000
rect 8200 3200 8500 4000
rect 10200 7000 10500 7100
rect 10200 4000 10300 7000
rect 10400 4000 10500 7000
rect 8800 3850 9200 3900
rect 8800 3650 8850 3850
rect 9150 3650 9200 3850
rect 8800 3600 9200 3650
rect 10200 3650 10500 4000
rect 10200 3450 10250 3650
rect 10450 3450 10500 3650
rect 10200 3200 10500 3450
rect 12200 7000 12500 7100
rect 12200 4000 12300 7000
rect 12400 4000 12500 7000
rect 12200 3200 12500 4000
rect -700 3100 17400 3200
rect -700 100 -400 3100
rect -300 100 1600 3100
rect 1700 100 3600 3100
rect 3700 100 5600 3100
rect 5700 100 8300 3100
rect 8400 100 11000 3100
rect 11100 100 13000 3100
rect 13100 100 15000 3100
rect 15100 100 17000 3100
rect 17100 100 17400 3100
rect -700 0 17400 100
<< via1 >>
rect 7550 7450 7850 7650
rect 8850 3650 9150 3850
<< metal2 >>
rect 7500 7650 7900 11200
rect 7500 7450 7550 7650
rect 7850 7450 7900 7650
rect 7500 7400 7900 7450
rect 8800 3850 9200 11200
rect 8800 3650 8850 3850
rect 9150 3650 9200 3850
rect 8800 3600 9200 3650
<< labels >>
flabel metal2 7700 11200 7700 11200 0 FreeSans 800 0 0 0 VBP
port 1 nsew
flabel metal2 9000 11200 9000 11200 0 FreeSans 800 0 0 0 VBN
port 2 nsew
flabel metal1 -700 1600 -700 1600 0 FreeSans 800 0 0 0 GND
port 4 nsew
flabel metal1 -700 9400 -700 9400 0 FreeSans 800 0 0 0 VDD
port 3 nsew
<< end >>

** sch_path: /home/lxbtlr/DTILO/schemas/inv_testbench.sch
**.subckt inv_testbench vout
*.opin vout
x1 net1 q0 vout n_inv
x2 net1 q1 q0 n_inv
x3 net1 q2 q1 n_inv
x4 net1 q3 q2 n_inv
x5 net1 vout q3 n_inv
V1 VDD GND 1.8
I1 VDD net2 {i_s}
XM1 VDD net2 net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 GND net2 net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.option wnflag=1
.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt


.param W=1 L=.15 i_s=.10n
.tran 1n 2n
.control
run
plot v(vout) v(q0) v(q1) v(q2) v(q3)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/lxbtlr/DTILO/schemas/n_inv.sym # of pins=3
** sym_path: /home/lxbtlr/DTILO/schemas/n_inv.sym
** sch_path: /home/lxbtlr/DTILO/schemas/n_inv.sch
.subckt n_inv VP Q A
*.ipin A
*.ipin VP
*.opin Q
XM1 Q A GND GND sky130_fd_pr__nfet_01v8 L={L} W={W} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Q A VP VDD sky130_fd_pr__pfet_01v8 L={L} W={W} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends

.GLOBAL VDD
.GLOBAL GND
.end

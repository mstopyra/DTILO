magic
tech sky130A
timestamp 1702655834
<< nwell >>
rect -7450 22050 -900 22100
rect -7450 22000 -6750 22050
rect -7450 18800 -6450 22000
rect -3850 21900 -1300 22050
rect -3900 20900 -1300 21900
rect -4000 19950 -1300 20900
rect 30000 21000 30200 21700
rect -4000 19750 100 19950
rect -7450 18700 -7150 18800
rect -6500 18700 -6450 18800
rect -3900 18700 -1300 19750
rect 30000 18850 30250 21000
rect 30000 15000 30200 18850
rect 36600 14950 37000 15300
<< pmos >>
rect -7150 18800 -6750 22000
<< pdiff >>
rect -7450 21900 -7150 22000
rect -7450 18900 -7350 21900
rect -7250 18900 -7150 21900
rect -7450 18800 -7150 18900
rect -6750 21900 -6450 22000
rect -6750 18900 -6650 21900
rect -6550 18900 -6450 21900
rect -6750 18800 -6450 18900
<< pdiffc >>
rect -7350 18900 -7250 21900
rect -6650 18900 -6550 21900
<< poly >>
rect -7150 22050 -900 22150
rect -7150 22000 -6750 22050
rect -7150 18750 -6750 18800
rect -4600 14550 -4450 22050
rect -4600 14400 -1000 14550
rect -4150 7150 -3800 7200
rect -4150 6950 -4100 7150
rect -3850 6950 -3800 7150
rect -4150 6900 -3800 6950
rect -3900 6750 -3800 6900
rect -3900 6700 -2950 6750
rect -3900 6650 -3050 6700
rect -3000 6650 -2950 6700
rect -3100 6600 -2950 6650
<< polycont >>
rect -4100 6950 -3850 7150
rect -3050 6650 -3000 6700
<< locali >>
rect -7550 18900 -7350 21900
rect -7250 18900 -7150 21900
rect -6750 18900 -6650 21900
rect -6550 18900 -6450 21900
rect -7350 18800 -7250 18900
rect -6650 15050 -6550 18900
rect 37020 16780 37210 16830
rect -6650 14950 -3700 15050
rect -3800 10100 -3700 14950
rect 36600 14900 36750 14950
rect 37020 14800 37070 16780
rect 40975 16330 40980 16350
rect 40935 16185 41085 16210
rect 40935 15770 40955 16185
rect 41855 16170 42140 16215
rect 36950 14750 37070 14800
rect 37170 15720 37260 15770
rect 40820 15750 40955 15770
rect -14050 10000 -3700 10100
rect -3200 14650 -2850 14750
rect 29950 14650 30050 14700
rect -14050 9550 -13950 10000
rect -4150 7150 -3800 7200
rect -4150 6950 -4100 7150
rect -3850 6950 -3800 7150
rect -3200 6950 -3100 14650
rect 3900 14500 11350 14600
rect 29950 14550 30150 14650
rect 37170 14630 37200 15720
rect 40820 14830 40850 15750
rect 40820 14805 41090 14830
rect 40820 14630 40850 14805
rect 42280 14790 42565 14835
rect 37170 14600 40850 14630
rect 30300 14550 30450 14600
rect 11250 13050 11350 14500
rect 30050 14450 30450 14550
rect 11250 12950 12400 13050
rect 12150 12750 12400 12950
rect 22950 12950 23200 13050
rect 22950 12750 23900 12950
rect 23700 11550 23900 12750
rect 30300 11550 30450 14450
rect 40820 13470 40850 14600
rect 40820 13445 41080 13470
rect 42685 13430 42835 13475
rect -4150 6900 -3800 6950
rect -3350 6800 -3050 6900
rect -3350 6550 -3250 6800
rect -3100 6700 -2950 6750
rect -3100 6650 -3050 6700
rect -3000 6650 -2950 6700
rect -3100 6600 -2950 6650
rect -4150 6450 -3250 6550
rect -4150 4400 -4050 6450
rect -4150 4100 -3800 4400
<< viali >>
rect -14850 9800 -14650 9900
<< metal1 >>
rect -7450 18800 -6450 22000
rect -4000 19950 -1300 20900
rect -4000 19750 100 19950
rect 7150 19750 12250 19950
rect 30000 18850 30250 21000
rect 36600 18850 36700 18900
rect -7450 14800 -7250 18800
rect -3350 15750 -1150 16050
rect 9150 15150 9250 17200
rect 36650 16280 36700 18850
rect 40850 16740 41055 16775
rect 41865 16740 42035 16775
rect 40850 16370 40895 16740
rect 40800 16335 40895 16370
rect 36650 16220 37020 16280
rect 37070 16220 37300 16280
rect 9150 15050 11200 15150
rect 36650 15100 36700 16220
rect 40985 15560 41065 15780
rect 40800 15480 41065 15560
rect 40800 15370 40895 15480
rect 41985 15380 42035 16740
rect 37130 15280 37220 15340
rect 36650 15050 36750 15100
rect -7450 14600 -3850 14800
rect -4050 14500 -3850 14600
rect -4050 14300 -3550 14500
rect -3700 14250 -3550 14300
rect -3700 14000 -2950 14250
rect -3700 10250 -3550 14000
rect 11100 10450 11200 15050
rect 36700 14950 36750 15050
rect 37130 14780 37190 15280
rect 40740 15275 40895 15370
rect 42300 15360 42485 15395
rect 36700 14550 36750 14750
rect 37000 14730 37190 14780
rect 36600 14500 36750 14550
rect 12100 13050 12450 13100
rect 12100 12750 12150 13050
rect 12400 12750 12450 13050
rect 12100 12700 12450 12750
rect 22900 13050 23250 13100
rect 22900 12750 22950 13050
rect 23200 12750 23250 13050
rect 22900 12700 23250 12750
rect 36600 13035 36650 14500
rect 40800 14400 40895 15275
rect 40750 14300 41070 14400
rect 42435 14030 42485 15360
rect 36600 12940 41045 13035
rect 36600 10700 36650 12940
rect 11000 10350 11200 10450
rect -14900 10100 -3550 10250
rect -14900 9900 -14600 10100
rect -14900 9800 -14850 9900
rect -14650 9800 -14600 9900
rect -14900 9750 -14600 9800
rect 21800 9300 24500 9650
rect 11000 7450 12150 7650
rect 21800 7500 22050 9300
rect -4200 7200 -3750 7250
rect -4200 6900 -4150 7200
rect -3800 6900 -3750 7200
rect -4200 6850 -3750 6900
rect -3600 5500 12350 6000
rect -4200 4400 -3750 4450
rect -4200 4100 -4150 4400
rect -3800 4100 -3750 4400
rect -4200 4050 -3750 4100
rect -3600 3950 -3050 5500
rect -4700 3400 -3050 3950
rect -4700 -1700 -4200 3400
rect -7250 -2200 -4200 -1700
<< via1 >>
rect 12150 12750 12400 13050
rect 22950 12750 23200 13050
rect -4150 6900 -3800 7200
rect -4150 4100 -3800 4400
<< metal2 >>
rect -12450 22200 11600 22300
rect 11500 11050 11600 22200
rect 22900 13050 23250 13100
rect 22900 12750 22950 13050
rect 23200 12750 23250 13050
rect 22900 12700 23250 12750
rect 11500 10950 12150 11050
use 4BIT_DAC_block  4BIT_DAC_block_0
timestamp 1702609360
transform 1 0 -18650 0 1 -8050
box 2000 -100 14900 18000
use BIASGEN_VBP_VBN  BIASGEN_VBP_VBN_0
timestamp 1701138250
transform 1 0 -21250 0 1 11000
box -700 -300 17400 11200
use f_div_four  f_div_four_0
timestamp 1702607528
transform 1 0 41030 0 1 12830
box -65 0 1735 1265
use f_div_three  f_div_three_0
timestamp 1702607100
transform 1 0 41040 0 1 14190
box -70 0 1320 1255
use f_div_two  f_div_two_0
timestamp 1702655834
transform 1 0 41035 0 1 15570
box -60 0 900 1255
use first_current_mirror  first_current_mirror_0
timestamp 1702612971
transform 1 0 13350 0 1 500
box -1250 -450 9550 21550
use FVF  FVF_0
timestamp 1702260771
transform 1 0 -2450 0 1 11100
box -650 -4450 13550 3400
use IN_AMP  IN_AMP_0
timestamp 1702573795
transform 1 0 30600 0 1 18350
box -400 -10450 6050 3350
use IN_AMP  IN_AMP_1
timestamp 1702573795
transform 1 0 24000 0 1 18350
box -400 -10450 6050 3350
use OUT_MIRROR  OUT_MIRROR_0
timestamp 1702603859
transform -1 0 36829 0 1 14705
box -175 -55 145 610
use RING_OSC  RING_OSC_0
timestamp 1702605233
transform 1 0 37210 0 1 14655
box -10 -5 3615 2235
use VCN_BIAS  VCN_BIAS_0
timestamp 1702585456
transform 1 0 -4000 0 1 20700
box 600 -6050 13150 1350
<< labels >>
flabel locali 42140 16190 42140 16190 0 FreeSans 800 0 0 0 Fdiv2
port 0 nsew
flabel locali 42565 14810 42565 14810 0 FreeSans 800 0 0 0 Fdiv3
port 4 nsew
flabel locali 42835 13450 42835 13450 0 FreeSans 800 0 0 0 Fdiv4
port 6 nsew
<< end >>

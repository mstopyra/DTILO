magic
tech sky130A
timestamp 1702585456
<< nwell >>
rect 2600 -2150 11150 1350
<< nmos >>
rect 1250 -5700 1650 -2500
rect 1950 -5700 2350 -2500
rect 3300 -5700 3700 -2500
rect 4000 -5700 4400 -2500
rect 5350 -5700 5750 -2500
rect 6050 -5700 6450 -2500
rect 7300 -5700 7700 -2500
rect 8000 -5700 8400 -2500
rect 9350 -5700 9750 -2500
rect 10050 -5700 10450 -2500
rect 11400 -5700 11800 -2500
rect 12100 -5700 12500 -2500
<< pmos >>
rect 2950 -2050 3350 1150
rect 4200 -2050 4600 1150
rect 4650 -2050 5050 1150
rect 5100 -2050 5500 1150
rect 5550 -2050 5950 1150
rect 6000 -2050 6400 1150
rect 7350 -2050 7750 1150
rect 7800 -2050 8200 1150
rect 8250 -2050 8650 1150
rect 8700 -2050 9100 1150
rect 9150 -2050 9550 1150
rect 10400 -2050 10800 1150
<< ndiff >>
rect 950 -2600 1250 -2500
rect 950 -5600 1050 -2600
rect 1150 -5600 1250 -2600
rect 950 -5700 1250 -5600
rect 1650 -2600 1950 -2500
rect 1650 -5600 1750 -2600
rect 1850 -5600 1950 -2600
rect 1650 -5700 1950 -5600
rect 2350 -2600 2650 -2500
rect 2350 -5600 2450 -2600
rect 2550 -5600 2650 -2600
rect 2350 -5700 2650 -5600
rect 3000 -2600 3300 -2500
rect 3000 -5600 3100 -2600
rect 3200 -5600 3300 -2600
rect 3000 -5700 3300 -5600
rect 3700 -2600 4000 -2500
rect 3700 -5600 3800 -2600
rect 3900 -5600 4000 -2600
rect 3700 -5700 4000 -5600
rect 4400 -2600 4700 -2500
rect 4400 -5600 4500 -2600
rect 4600 -5600 4700 -2600
rect 4400 -5700 4700 -5600
rect 5050 -2600 5350 -2500
rect 5050 -5600 5150 -2600
rect 5250 -5600 5350 -2600
rect 5050 -5700 5350 -5600
rect 5750 -2600 6050 -2500
rect 5750 -5600 5850 -2600
rect 5950 -5600 6050 -2600
rect 5750 -5650 6050 -5600
rect 5750 -5700 5800 -5650
rect 5900 -5700 6050 -5650
rect 6450 -2600 6750 -2500
rect 7000 -2600 7300 -2500
rect 6450 -5600 6550 -2600
rect 6650 -5600 6750 -2600
rect 7000 -5600 7100 -2600
rect 7200 -5600 7300 -2600
rect 6450 -5700 6750 -5600
rect 7000 -5700 7300 -5600
rect 7700 -2600 8000 -2500
rect 7700 -5600 7800 -2600
rect 7900 -5600 8000 -2600
rect 7700 -5650 8000 -5600
rect 7700 -5700 7850 -5650
rect 7950 -5700 8000 -5650
rect 8400 -2600 8700 -2500
rect 8400 -5600 8500 -2600
rect 8600 -5600 8700 -2600
rect 8400 -5700 8700 -5600
rect 9050 -2600 9350 -2500
rect 9050 -5600 9150 -2600
rect 9250 -5600 9350 -2600
rect 9050 -5700 9350 -5600
rect 9750 -2600 10050 -2500
rect 9750 -5600 9850 -2600
rect 9950 -5600 10050 -2600
rect 9750 -5700 10050 -5600
rect 10450 -2600 10750 -2500
rect 10450 -5600 10550 -2600
rect 10650 -5600 10750 -2600
rect 10450 -5700 10750 -5600
rect 11100 -2600 11400 -2500
rect 11100 -5600 11200 -2600
rect 11300 -5600 11400 -2600
rect 11100 -5700 11400 -5600
rect 11800 -2600 12100 -2500
rect 11800 -5600 11900 -2600
rect 12000 -5600 12100 -2600
rect 11800 -5700 12100 -5600
rect 12500 -2600 12800 -2500
rect 12500 -5600 12600 -2600
rect 12700 -5600 12800 -2600
rect 12500 -5700 12800 -5600
<< pdiff >>
rect 2650 1050 2950 1150
rect 2650 -1950 2750 1050
rect 2850 -1950 2950 1050
rect 2650 -2050 2950 -1950
rect 3350 1050 3650 1150
rect 3900 1050 4200 1150
rect 3350 -1950 3450 1050
rect 3550 -1950 3650 1050
rect 3900 -1950 4000 1050
rect 4100 -1950 4200 1050
rect 3350 -2050 3650 -1950
rect 3900 -2050 4200 -1950
rect 4600 -2050 4650 1150
rect 5050 -2050 5100 1150
rect 5500 -2050 5550 1150
rect 5950 -2050 6000 1150
rect 6400 1050 6700 1150
rect 6400 -1950 6500 1050
rect 6600 -1950 6700 1050
rect 6400 -2050 6700 -1950
rect 7050 1050 7350 1150
rect 7050 -1950 7150 1050
rect 7250 -1950 7350 1050
rect 7050 -2050 7350 -1950
rect 7750 -2050 7800 1150
rect 8200 -2050 8250 1150
rect 8650 -2050 8700 1150
rect 9100 -2050 9150 1150
rect 9550 1050 9850 1150
rect 10100 1050 10400 1150
rect 9550 -1950 9650 1050
rect 9750 -1950 9850 1050
rect 10100 -1950 10200 1050
rect 10300 -1950 10400 1050
rect 9550 -2050 9850 -1950
rect 10100 -2050 10400 -1950
rect 10800 1050 11100 1150
rect 10800 -1950 10900 1050
rect 11000 -1950 11100 1050
rect 10800 -2050 11100 -1950
<< ndiffc >>
rect 1050 -5600 1150 -2600
rect 1750 -5600 1850 -2600
rect 2450 -5600 2550 -2600
rect 3100 -5600 3200 -2600
rect 3800 -5600 3900 -2600
rect 4500 -5600 4600 -2600
rect 5150 -5600 5250 -2600
rect 5850 -5600 5950 -2600
rect 6550 -5600 6650 -2600
rect 7100 -5600 7200 -2600
rect 7800 -5600 7900 -2600
rect 8500 -5600 8600 -2600
rect 9150 -5600 9250 -2600
rect 9850 -5600 9950 -2600
rect 10550 -5600 10650 -2600
rect 11200 -5600 11300 -2600
rect 11900 -5600 12000 -2600
rect 12600 -5600 12700 -2600
<< pdiffc >>
rect 2750 -1950 2850 1050
rect 3450 -1950 3550 1050
rect 4000 -1950 4100 1050
rect 6500 -1950 6600 1050
rect 7150 -1950 7250 1050
rect 9650 -1950 9750 1050
rect 10200 -1950 10300 1050
rect 10900 -1950 11000 1050
<< psubdiff >>
rect 650 -2600 900 -2500
rect 650 -5600 750 -2600
rect 800 -5600 900 -2600
rect 650 -5700 900 -5600
rect 2700 -2600 2950 -2500
rect 2700 -5600 2800 -2600
rect 2850 -5600 2950 -2600
rect 2700 -5700 2950 -5600
rect 4750 -2600 5000 -2500
rect 4750 -5600 4850 -2600
rect 4900 -5600 5000 -2600
rect 4750 -5700 5000 -5600
rect 6750 -2600 7000 -2500
rect 6750 -5600 6850 -2600
rect 6900 -5600 7000 -2600
rect 6750 -5700 7000 -5600
rect 8750 -2600 9000 -2500
rect 8750 -5600 8850 -2600
rect 8900 -5600 9000 -2600
rect 8750 -5700 9000 -5600
rect 10800 -2600 11050 -2500
rect 10800 -5600 10900 -2600
rect 10950 -5600 11050 -2600
rect 10800 -5700 11050 -5600
rect 12850 -2600 13100 -2500
rect 12850 -5600 12950 -2600
rect 13000 -5600 13100 -2600
rect 12850 -5700 13100 -5600
<< nsubdiff >>
rect 3650 1050 3900 1150
rect 3650 -1950 3750 1050
rect 3800 -1950 3900 1050
rect 3650 -2050 3900 -1950
rect 6750 1050 7000 1150
rect 6750 -1950 6850 1050
rect 6900 -1950 7000 1050
rect 6750 -2050 7000 -1950
rect 9850 1050 10100 1150
rect 9850 -1950 9950 1050
rect 10000 -1950 10100 1050
rect 9850 -2050 10100 -1950
<< psubdiffcont >>
rect 750 -5600 800 -2600
rect 2800 -5600 2850 -2600
rect 4850 -5600 4900 -2600
rect 6850 -5600 6900 -2600
rect 8850 -5600 8900 -2600
rect 10900 -5600 10950 -2600
rect 12950 -5600 13000 -2600
<< nsubdiffcont >>
rect 3750 -1950 3800 1050
rect 6850 -1950 6900 1050
rect 9950 -1950 10000 1050
<< poly >>
rect 2950 1300 3100 1350
rect 2950 1250 3000 1300
rect 3050 1250 6400 1300
rect 2950 1200 6400 1250
rect 2950 1150 3350 1200
rect 4200 1150 4600 1200
rect 4650 1150 5050 1200
rect 5100 1150 5500 1200
rect 5550 1150 5950 1200
rect 6000 1150 6400 1200
rect 7350 1200 10800 1300
rect 7350 1150 7750 1200
rect 7800 1150 8200 1200
rect 8250 1150 8650 1200
rect 8700 1150 9100 1200
rect 9150 1150 9550 1200
rect 10400 1150 10800 1200
rect 2950 -2100 3350 -2050
rect 4200 -2100 4600 -2050
rect 4650 -2100 5050 -2050
rect 5100 -2100 5500 -2050
rect 5550 -2100 5950 -2050
rect 6000 -2100 6400 -2050
rect 7350 -2100 7750 -2050
rect 7800 -2100 8200 -2050
rect 8250 -2100 8650 -2050
rect 8700 -2100 9100 -2050
rect 9150 -2100 9550 -2050
rect 10400 -2100 10800 -2050
rect 1250 -2350 1400 -2300
rect 2450 -2350 2600 -2300
rect 3050 -2350 3200 -2300
rect 3750 -2350 3900 -2300
rect 4450 -2350 4600 -2300
rect 5100 -2350 5250 -2300
rect 6500 -2350 6650 -2300
rect 7100 -2350 7250 -2300
rect 8500 -2350 8650 -2300
rect 9150 -2350 9300 -2300
rect 9850 -2350 10000 -2300
rect 10550 -2350 10700 -2300
rect 11150 -2350 11300 -2300
rect 12350 -2350 12500 -2300
rect 1250 -2400 1300 -2350
rect 1350 -2400 2500 -2350
rect 2550 -2400 3100 -2350
rect 3150 -2400 3800 -2350
rect 3850 -2400 4500 -2350
rect 4550 -2400 5150 -2350
rect 5200 -2400 6550 -2350
rect 6600 -2400 7150 -2350
rect 7200 -2400 8550 -2350
rect 8600 -2400 9200 -2350
rect 9250 -2400 9900 -2350
rect 9950 -2400 10600 -2350
rect 10650 -2400 11200 -2350
rect 11250 -2400 12400 -2350
rect 12450 -2400 12500 -2350
rect 1250 -2450 12500 -2400
rect 1250 -2500 1650 -2450
rect 1950 -2500 2350 -2450
rect 3300 -2500 3700 -2450
rect 4000 -2500 4400 -2450
rect 5350 -2500 5750 -2450
rect 6050 -2500 6450 -2450
rect 7300 -2500 7700 -2450
rect 8000 -2500 8400 -2450
rect 9350 -2500 9750 -2450
rect 10050 -2500 10450 -2450
rect 11400 -2500 11800 -2450
rect 12100 -2500 12500 -2450
rect 1250 -5750 1650 -5700
rect 1950 -5750 2350 -5700
rect 3300 -5750 3700 -5700
rect 4000 -5750 4400 -5700
rect 5350 -5750 5750 -5700
rect 6050 -5750 6450 -5700
rect 7300 -5750 7700 -5700
rect 8000 -5750 8400 -5700
rect 9350 -5750 9750 -5700
rect 10050 -5750 10450 -5700
rect 11400 -5750 11800 -5700
rect 12100 -5750 12500 -5700
<< polycont >>
rect 3000 1250 3050 1300
rect 1300 -2400 1350 -2350
rect 2500 -2400 2550 -2350
rect 3100 -2400 3150 -2350
rect 3800 -2400 3850 -2350
rect 4500 -2400 4550 -2350
rect 5150 -2400 5200 -2350
rect 6550 -2400 6600 -2350
rect 7150 -2400 7200 -2350
rect 8550 -2400 8600 -2350
rect 9200 -2400 9250 -2350
rect 9900 -2400 9950 -2350
rect 10600 -2400 10650 -2350
rect 11200 -2400 11250 -2350
rect 12400 -2400 12450 -2350
<< locali >>
rect 2600 1300 3100 1350
rect 2600 1250 3000 1300
rect 3050 1250 3100 1300
rect 2600 1200 3100 1250
rect 2700 1050 2900 1100
rect 2700 -1850 2750 1050
rect 1250 -1950 2750 -1850
rect 2850 -1950 2900 1050
rect 1250 -2000 2900 -1950
rect 3400 1050 4150 1100
rect 3400 -1950 3450 1050
rect 3550 -1950 3750 1050
rect 3800 -1950 4000 1050
rect 4100 -1950 4150 1050
rect 3400 -2000 4150 -1950
rect 6450 1050 6650 1100
rect 6450 -1950 6500 1050
rect 6600 -1950 6650 1050
rect 6450 -2000 6650 -1950
rect 6800 1050 6950 1100
rect 6800 -1950 6850 1050
rect 6900 -1950 6950 1050
rect 6800 -2000 6950 -1950
rect 7100 1050 7300 1100
rect 7100 -1950 7150 1050
rect 7250 -1950 7300 1050
rect 7100 -2000 7300 -1950
rect 9600 1050 10350 1100
rect 9600 -1950 9650 1050
rect 9750 -1950 9950 1050
rect 10000 -1950 10200 1050
rect 10300 -1950 10350 1050
rect 9600 -2000 10350 -1950
rect 10850 1050 11050 1100
rect 10850 -1950 10900 1050
rect 11000 -1850 11050 1050
rect 11000 -1950 12500 -1850
rect 10850 -2000 12500 -1950
rect 1250 -2350 1400 -2000
rect 6500 -2100 6650 -2000
rect 7100 -2100 7250 -2000
rect 6500 -2200 7250 -2100
rect 1250 -2400 1300 -2350
rect 1350 -2400 1400 -2350
rect 1250 -2450 1400 -2400
rect 2450 -2350 2600 -2300
rect 2450 -2400 2500 -2350
rect 2550 -2400 2600 -2350
rect 2450 -2550 2600 -2400
rect 3050 -2350 3200 -2300
rect 3050 -2400 3100 -2350
rect 3150 -2400 3200 -2350
rect 3050 -2550 3200 -2400
rect 3750 -2350 3900 -2300
rect 3750 -2400 3800 -2350
rect 3850 -2400 3900 -2350
rect 3750 -2550 3900 -2400
rect 4450 -2350 4600 -2300
rect 4450 -2400 4500 -2350
rect 4550 -2400 4600 -2350
rect 4450 -2550 4600 -2400
rect 5100 -2350 5250 -2300
rect 5100 -2400 5150 -2350
rect 5200 -2400 5250 -2350
rect 5100 -2550 5250 -2400
rect 6500 -2350 6650 -2200
rect 6500 -2400 6550 -2350
rect 6600 -2400 6650 -2350
rect 6500 -2550 6650 -2400
rect 7100 -2350 7250 -2200
rect 7100 -2400 7150 -2350
rect 7200 -2400 7250 -2350
rect 7100 -2550 7250 -2400
rect 8500 -2350 8650 -2300
rect 8500 -2400 8550 -2350
rect 8600 -2400 8650 -2350
rect 8500 -2550 8650 -2400
rect 9150 -2350 9300 -2300
rect 9150 -2400 9200 -2350
rect 9250 -2400 9300 -2350
rect 9150 -2550 9300 -2400
rect 9850 -2350 10000 -2300
rect 9850 -2400 9900 -2350
rect 9950 -2400 10000 -2350
rect 9850 -2550 10000 -2400
rect 10550 -2350 10700 -2300
rect 10550 -2400 10600 -2350
rect 10650 -2400 10700 -2350
rect 10550 -2550 10700 -2400
rect 11150 -2350 11300 -2300
rect 11150 -2400 11200 -2350
rect 11250 -2400 11300 -2350
rect 11150 -2550 11300 -2400
rect 12350 -2350 12500 -2000
rect 12350 -2400 12400 -2350
rect 12450 -2400 12500 -2350
rect 12350 -2450 12500 -2400
rect 700 -2600 850 -2550
rect 700 -5600 750 -2600
rect 800 -5600 850 -2600
rect 700 -5650 850 -5600
rect 1000 -2600 1200 -2550
rect 1000 -5600 1050 -2600
rect 1150 -5600 1200 -2600
rect 1000 -5650 1200 -5600
rect 1700 -2600 1900 -2550
rect 1700 -5600 1750 -2600
rect 1850 -5600 1900 -2600
rect 1700 -5650 1900 -5600
rect 2400 -2600 2600 -2550
rect 2400 -5600 2450 -2600
rect 2550 -5600 2600 -2600
rect 2400 -5650 2600 -5600
rect 2750 -2600 2900 -2550
rect 2750 -5600 2800 -2600
rect 2850 -5600 2900 -2600
rect 2750 -5650 2900 -5600
rect 3050 -2600 3250 -2550
rect 3050 -5600 3100 -2600
rect 3200 -5600 3250 -2600
rect 3050 -5650 3250 -5600
rect 3750 -2600 3950 -2550
rect 3750 -5600 3800 -2600
rect 3900 -5600 3950 -2600
rect 3750 -5650 3950 -5600
rect 4450 -2600 4650 -2550
rect 4450 -5600 4500 -2600
rect 4600 -5600 4650 -2600
rect 4450 -5650 4650 -5600
rect 4800 -2600 4950 -2550
rect 4800 -5600 4850 -2600
rect 4900 -5600 4950 -2600
rect 4800 -5650 4950 -5600
rect 5100 -2600 5300 -2550
rect 5100 -5600 5150 -2600
rect 5250 -5600 5300 -2600
rect 5100 -5650 5300 -5600
rect 5800 -2600 6000 -2550
rect 5800 -5600 5850 -2600
rect 5950 -5600 6000 -2600
rect 5800 -5650 6000 -5600
rect 6500 -2600 7250 -2550
rect 6500 -5600 6550 -2600
rect 6650 -5600 6850 -2600
rect 6900 -5600 7100 -2600
rect 7200 -5600 7250 -2600
rect 6500 -5650 7250 -5600
rect 7750 -2600 7950 -2550
rect 7750 -5600 7800 -2600
rect 7900 -5600 7950 -2600
rect 7750 -5650 7950 -5600
rect 8450 -2600 8650 -2550
rect 8450 -5600 8500 -2600
rect 8600 -5600 8650 -2600
rect 8450 -5650 8650 -5600
rect 8800 -2600 8950 -2550
rect 8800 -5600 8850 -2600
rect 8900 -5600 8950 -2600
rect 8800 -5650 8950 -5600
rect 9100 -2600 9300 -2550
rect 9100 -5600 9150 -2600
rect 9250 -5600 9300 -2600
rect 9100 -5650 9300 -5600
rect 9800 -2600 10000 -2550
rect 9800 -5600 9850 -2600
rect 9950 -5600 10000 -2600
rect 9800 -5650 10000 -5600
rect 10500 -2600 10700 -2550
rect 10500 -5600 10550 -2600
rect 10650 -5600 10700 -2600
rect 10500 -5650 10700 -5600
rect 10850 -2600 11000 -2550
rect 10850 -5600 10900 -2600
rect 10950 -5600 11000 -2600
rect 10850 -5650 11000 -5600
rect 11150 -2600 11350 -2550
rect 11150 -5600 11200 -2600
rect 11300 -5600 11350 -2600
rect 11150 -5650 11350 -5600
rect 11850 -2600 12050 -2550
rect 11850 -5600 11900 -2600
rect 12000 -5600 12050 -2600
rect 11850 -5650 12050 -5600
rect 12550 -2600 12750 -2550
rect 12550 -5600 12600 -2600
rect 12700 -5600 12750 -2600
rect 12550 -5650 12750 -5600
rect 12900 -2600 13050 -2550
rect 12900 -5600 12950 -2600
rect 13000 -5600 13050 -2600
rect 12900 -5650 13050 -5600
rect 1100 -5950 1200 -5650
rect 1800 -5800 1900 -5650
rect 5800 -5800 5900 -5650
rect 7850 -5800 7950 -5650
rect 11850 -5800 11950 -5650
rect 1800 -5900 11950 -5800
rect 12550 -5950 12650 -5650
rect 13050 -5950 13150 -5800
rect 1100 -6050 13150 -5950
<< viali >>
rect 3750 -900 3800 150
rect 6850 -900 6900 150
rect 9950 -900 10000 150
rect 750 -4600 800 -3550
rect 2800 -4600 2850 -3550
rect 4850 -4600 4900 -3550
rect 6550 -4600 6650 -3550
rect 6850 -4600 6900 -3550
rect 7100 -4600 7200 -3550
rect 8850 -4600 8900 -3550
rect 10900 -4600 10950 -3550
rect 12950 -4600 13000 -3550
<< metal1 >>
rect 2600 150 11150 200
rect 2600 -900 3750 150
rect 3800 -900 6850 150
rect 6900 -900 9950 150
rect 10000 -900 11150 150
rect 2600 -950 11150 -900
rect 600 -3550 13150 -3500
rect 600 -4600 750 -3550
rect 800 -4600 2800 -3550
rect 2850 -4600 4850 -3550
rect 4900 -4600 6550 -3550
rect 6650 -4600 6850 -3550
rect 6900 -4600 7100 -3550
rect 7200 -4600 8850 -3550
rect 8900 -4600 10900 -3550
rect 10950 -4600 12950 -3550
rect 13000 -4600 13150 -3550
rect 600 -4650 13150 -4600
<< labels >>
flabel locali 13150 -5950 13150 -5950 0 FreeSans 800 0 0 0 VCN
port 1 nsew
flabel metal1 600 -4000 600 -4000 0 FreeSans 800 0 0 0 GND
port 2 nsew
flabel metal1 2600 -400 2600 -400 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel locali 2600 1250 2600 1250 0 FreeSans 800 0 0 0 VG
port 4 nsew
<< end >>

magic
tech sky130A
timestamp 1702603859
<< nwell >>
rect -175 290 -20 575
rect -175 135 145 290
<< nmos >>
rect -105 0 -90 100
rect 60 0 75 100
<< pmos >>
rect -105 155 -90 555
rect 60 155 75 255
<< ndiff >>
rect -155 85 -105 100
rect -155 15 -140 85
rect -120 15 -105 85
rect -155 0 -105 15
rect -90 85 -40 100
rect 10 85 60 100
rect -90 15 -75 85
rect -55 15 -40 85
rect 10 15 25 85
rect 45 15 60 85
rect -90 0 -40 15
rect 10 0 60 15
rect 75 85 125 100
rect 75 15 90 85
rect 110 15 125 85
rect 75 0 125 15
<< pdiff >>
rect -155 240 -105 555
rect -155 170 -140 240
rect -120 170 -105 240
rect -155 155 -105 170
rect -90 255 -55 555
rect -90 240 -40 255
rect 10 240 60 255
rect -90 170 -75 240
rect -55 170 -40 240
rect 10 170 25 240
rect 45 170 60 240
rect -90 155 -40 170
rect 10 155 60 170
rect 75 240 125 255
rect 75 170 90 240
rect 110 170 125 240
rect 75 155 125 170
<< ndiffc >>
rect -140 15 -120 85
rect -75 15 -55 85
rect 25 15 45 85
rect 90 15 110 85
<< pdiffc >>
rect -140 170 -120 240
rect -75 170 -55 240
rect 25 170 45 240
rect 90 170 110 240
<< psubdiff >>
rect -40 85 10 100
rect -40 15 -25 85
rect -5 15 10 85
rect -40 0 10 15
<< nsubdiff >>
rect -40 240 10 255
rect -40 170 -25 240
rect -5 170 10 240
rect -40 155 10 170
<< psubdiffcont >>
rect -25 15 -5 85
<< nsubdiffcont >>
rect -25 170 -5 240
<< poly >>
rect -130 600 -90 610
rect -130 580 -120 600
rect -100 580 -90 600
rect -130 570 -30 580
rect -105 565 -30 570
rect -105 555 -90 565
rect -45 290 -30 565
rect -45 275 75 290
rect 60 255 75 275
rect -105 140 -90 155
rect 60 140 75 155
rect -105 100 -90 115
rect 60 100 75 115
rect -105 -15 -90 0
rect 60 -15 75 0
rect -105 -25 75 -15
rect -105 -45 -95 -25
rect -75 -30 75 -25
rect -75 -45 -65 -30
rect -105 -55 -65 -45
<< polycont >>
rect -120 580 -100 600
rect -95 -45 -75 -25
<< locali >>
rect -130 600 -90 610
rect -130 580 -120 600
rect -100 580 -90 600
rect -130 570 -90 580
rect -130 250 -110 570
rect -150 240 -110 250
rect -150 170 -140 240
rect -120 170 -110 240
rect -150 160 -110 170
rect -85 240 55 250
rect -85 170 -75 240
rect -55 170 -25 240
rect -5 170 25 240
rect 45 170 55 240
rect -85 160 55 170
rect 80 240 120 250
rect 80 170 90 240
rect 110 170 120 240
rect 80 160 120 170
rect -130 135 -110 160
rect -130 115 100 135
rect 80 95 100 115
rect -150 85 -110 95
rect -150 15 -140 85
rect -120 15 -110 85
rect -150 5 -110 15
rect -85 85 55 95
rect -85 15 -75 85
rect -55 15 -25 85
rect -5 15 25 85
rect 45 15 55 85
rect -85 5 55 15
rect 80 85 120 95
rect 80 15 90 85
rect 110 15 120 85
rect 80 5 120 15
rect -85 -15 -65 5
rect -105 -25 -65 -15
rect -105 -45 -95 -25
rect -75 -45 -65 -25
rect -105 -55 -65 -45
<< viali >>
rect -75 170 -55 240
rect -25 170 -5 240
rect 25 170 45 240
rect -75 15 -55 85
rect -25 15 -5 85
rect 25 15 45 85
<< metal1 >>
rect -175 240 145 255
rect -175 170 -75 240
rect -55 170 -25 240
rect -5 170 25 240
rect 45 170 145 240
rect -175 155 145 170
rect -175 85 145 100
rect -175 15 -75 85
rect -55 15 -25 85
rect -5 15 25 85
rect 45 15 145 85
rect -175 0 145 15
<< labels >>
flabel metal1 -175 45 -175 45 0 FreeSans 400 0 0 0 amp_i_out
port 0 nsew
flabel metal1 145 200 145 200 0 FreeSans 400 0 0 0 RO_in
port 1 nsew
flabel metal1 -175 205 -175 205 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 145 50 145 50 0 FreeSans 400 0 0 0 GND
port 3 nsew
<< end >>

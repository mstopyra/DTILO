magic
tech sky130A
timestamp 1702573795
<< nwell >>
rect -400 -3350 6000 3350
rect -200 -3400 -100 -3350
<< nmos >>
rect -50 -10250 350 -7050
rect 1250 -10250 1650 -3850
rect 1950 -10250 2350 -3850
rect 3250 -10250 3650 -3850
rect 3950 -10250 4350 -3850
rect 5250 -10250 5650 -3850
<< pmos >>
rect -50 -50 350 3150
rect 1250 -3250 1650 3150
rect 1950 -3250 2350 3150
rect 3250 -3250 3650 3150
rect 3950 -3250 4350 3150
rect 5250 -3250 5650 3150
<< ndiff >>
rect 600 -7050 650 -3850
rect 950 -3950 1250 -3850
rect -350 -7150 -50 -7050
rect -350 -10150 -250 -7150
rect -150 -10150 -50 -7150
rect -350 -10250 -50 -10150
rect 350 -7150 650 -7050
rect 350 -10150 450 -7150
rect 550 -10150 650 -7150
rect 950 -10150 1050 -3950
rect 1150 -10150 1250 -3950
rect 350 -10250 650 -10150
rect 950 -10250 1250 -10150
rect 1650 -3950 1950 -3850
rect 1650 -10150 1750 -3950
rect 1850 -10150 1950 -3950
rect 1650 -10250 1950 -10150
rect 2350 -3950 2650 -3850
rect 2950 -3950 3250 -3850
rect 2350 -10150 2450 -3950
rect 2550 -10150 2650 -3950
rect 2950 -10150 3050 -3950
rect 3150 -10150 3250 -3950
rect 2350 -10250 2650 -10150
rect 2950 -10250 3250 -10150
rect 3650 -3950 3950 -3850
rect 3650 -10150 3750 -3950
rect 3850 -10150 3950 -3950
rect 3650 -10250 3950 -10150
rect 4350 -3950 4650 -3850
rect 4950 -3950 5250 -3850
rect 4350 -10150 4450 -3950
rect 4550 -10150 4650 -3950
rect 4950 -10150 5050 -3950
rect 5150 -10150 5250 -3950
rect 4350 -10250 4650 -10150
rect 4950 -10250 5250 -10150
rect 5650 -3950 5950 -3850
rect 5650 -10150 5750 -3950
rect 5850 -10150 5950 -3950
rect 5650 -10250 5950 -10150
<< pdiff >>
rect -350 3050 -50 3150
rect -350 50 -250 3050
rect -150 50 -50 3050
rect -350 -50 -50 50
rect 350 3050 650 3150
rect 950 3050 1250 3150
rect 350 50 450 3050
rect 550 50 650 3050
rect 350 -50 650 50
rect 600 -3250 650 -50
rect 950 -3150 1050 3050
rect 1150 -3150 1250 3050
rect 950 -3250 1250 -3150
rect 1650 3050 1950 3150
rect 1650 -3150 1750 3050
rect 1850 -3150 1950 3050
rect 1650 -3250 1950 -3150
rect 2350 3050 2650 3150
rect 2950 3050 3250 3150
rect 2350 -3150 2450 3050
rect 2550 -3150 2650 3050
rect 2950 -3150 3050 3050
rect 3150 -3150 3250 3050
rect 2350 -3250 2650 -3150
rect 2950 -3250 3250 -3150
rect 3650 3050 3950 3150
rect 3650 -3150 3750 3050
rect 3850 -3150 3950 3050
rect 3650 -3250 3950 -3150
rect 4350 3050 4650 3150
rect 4950 3050 5250 3150
rect 4350 -3150 4450 3050
rect 4550 -3150 4650 3050
rect 4950 -3150 5050 3050
rect 5150 -3150 5250 3050
rect 4350 -3250 4650 -3150
rect 4950 -3250 5250 -3150
rect 5650 3050 5950 3150
rect 5650 -3150 5750 3050
rect 5850 -3150 5950 3050
rect 5650 -3250 5950 -3150
<< ndiffc >>
rect -250 -10150 -150 -7150
rect 450 -10150 550 -7150
rect 1050 -10150 1150 -3950
rect 1750 -10150 1850 -3950
rect 2450 -10150 2550 -3950
rect 3050 -10150 3150 -3950
rect 3750 -10150 3850 -3950
rect 4450 -10150 4550 -3950
rect 5050 -10150 5150 -3950
rect 5750 -10150 5850 -3950
<< pdiffc >>
rect -250 50 -150 3050
rect 450 50 550 3050
rect 1050 -3150 1150 3050
rect 1750 -3150 1850 3050
rect 2450 -3150 2550 3050
rect 3050 -3150 3150 3050
rect 3750 -3150 3850 3050
rect 4450 -3150 4550 3050
rect 5050 -3150 5150 3050
rect 5750 -3150 5850 3050
<< psubdiff >>
rect 650 -3950 950 -3850
rect 650 -10150 750 -3950
rect 850 -10150 950 -3950
rect 650 -10250 950 -10150
rect 2650 -3950 2950 -3850
rect 2650 -10150 2750 -3950
rect 2850 -10150 2950 -3950
rect 2650 -10250 2950 -10150
rect 4650 -3950 4950 -3850
rect 4650 -10150 4750 -3950
rect 4850 -10150 4950 -3950
rect 4650 -10250 4950 -10150
<< nsubdiff >>
rect 650 3050 950 3150
rect 650 -3150 750 3050
rect 850 -3150 950 3050
rect 650 -3250 950 -3150
rect 2650 3050 2950 3150
rect 2650 -3150 2750 3050
rect 2850 -3150 2950 3050
rect 2650 -3250 2950 -3150
rect 4650 3050 4950 3150
rect 4650 -3150 4750 3050
rect 4850 -3150 4950 3050
rect 4650 -3250 4950 -3150
<< psubdiffcont >>
rect 750 -10150 850 -3950
rect 2750 -10150 2850 -3950
rect 4750 -10150 4850 -3950
<< nsubdiffcont >>
rect 750 -3150 850 3050
rect 2750 -3150 2850 3050
rect 4750 -3150 4850 3050
<< poly >>
rect -50 3300 100 3350
rect -50 3250 0 3300
rect 50 3250 5650 3300
rect -50 3200 5650 3250
rect -50 3150 350 3200
rect 1250 3150 1650 3200
rect 1950 3150 2350 3200
rect 3250 3150 3650 3200
rect 3950 3150 4350 3200
rect 5250 3150 5650 3200
rect -50 -100 350 -50
rect 1250 -3300 1650 -3250
rect 1950 -3300 2350 -3250
rect 3250 -3300 3650 -3250
rect 3950 -3300 4350 -3250
rect 5250 -3300 5650 -3250
rect 1250 -3850 1650 -3800
rect 1950 -3850 2350 -3800
rect 3250 -3850 3650 -3800
rect 3950 -3850 4350 -3800
rect 5250 -3850 5650 -3800
rect -50 -7050 350 -7000
rect -50 -10300 350 -10250
rect 1250 -10300 1650 -10250
rect 1950 -10300 2350 -10250
rect 3250 -10300 3650 -10250
rect 3950 -10300 4350 -10250
rect 5250 -10300 5650 -10250
rect -50 -10350 5650 -10300
rect -50 -10400 0 -10350
rect 50 -10400 5650 -10350
rect -50 -10450 100 -10400
<< polycont >>
rect 0 3250 50 3300
rect 0 -10400 50 -10350
<< locali >>
rect -50 3300 100 3350
rect -200 3250 0 3300
rect 50 3250 100 3300
rect -200 3200 100 3250
rect -200 3100 -100 3200
rect -300 3050 -100 3100
rect -300 50 -250 3050
rect -150 50 -100 3050
rect -300 0 -100 50
rect 400 3050 1200 3100
rect 400 50 450 3050
rect 550 50 750 3050
rect 400 0 750 50
rect -200 -3600 -100 0
rect 700 -3150 750 0
rect 850 -3150 1050 3050
rect 1150 -3150 1200 3050
rect 700 -3200 1200 -3150
rect 1700 3050 1900 3100
rect 1700 -3150 1750 3050
rect 1850 -3150 1900 3050
rect 1700 -3200 1900 -3150
rect 2400 3050 3200 3100
rect 2400 -3150 2450 3050
rect 2550 -3150 2750 3050
rect 2850 -3150 3050 3050
rect 3150 -3150 3200 3050
rect 2400 -3200 3200 -3150
rect 3700 3050 3900 3100
rect 3700 -3150 3750 3050
rect 3850 -3150 3900 3050
rect 3700 -3200 3900 -3150
rect 4400 3050 5200 3100
rect 4400 -3150 4450 3050
rect 4550 -3150 4750 3050
rect 4850 -3150 5050 3050
rect 5150 -3150 5200 3050
rect 4400 -3200 5200 -3150
rect 5700 3050 5900 3100
rect 5700 -3150 5750 3050
rect 5850 -3150 5900 3050
rect 5700 -3200 5900 -3150
rect 1800 -3400 1900 -3200
rect 2650 -3250 2950 -3200
rect 3750 -3400 3850 -3200
rect 4650 -3250 4950 -3200
rect 5700 -3400 5800 -3200
rect 1800 -3500 6050 -3400
rect -200 -3700 5800 -3600
rect 5950 -3700 6050 -3500
rect 1800 -3900 1900 -3700
rect 2650 -3900 2950 -3850
rect 3750 -3900 3850 -3700
rect 4650 -3900 4950 -3850
rect 5700 -3900 5800 -3700
rect 700 -3950 1200 -3900
rect -300 -7150 -100 -6800
rect 700 -7100 750 -3950
rect -300 -10150 -250 -7150
rect -150 -10150 -100 -7150
rect -300 -10200 -100 -10150
rect 400 -7150 750 -7100
rect 400 -10150 450 -7150
rect 550 -10150 750 -7150
rect 850 -10150 1050 -3950
rect 1150 -10150 1200 -3950
rect 400 -10200 1200 -10150
rect 1700 -3950 1900 -3900
rect 1700 -10150 1750 -3950
rect 1850 -10150 1900 -3950
rect 1700 -10200 1900 -10150
rect 2400 -3950 3200 -3900
rect 2400 -10150 2450 -3950
rect 2550 -10150 2750 -3950
rect 2850 -10150 3050 -3950
rect 3150 -10150 3200 -3950
rect 2400 -10200 3200 -10150
rect 3700 -3950 3900 -3900
rect 3700 -10150 3750 -3950
rect 3850 -10150 3900 -3950
rect 3700 -10200 3900 -10150
rect 4400 -3950 5200 -3900
rect 4400 -10150 4450 -3950
rect 4550 -10150 4750 -3950
rect 4850 -10150 5050 -3950
rect 5150 -10150 5200 -3950
rect 4400 -10200 5200 -10150
rect 5700 -3950 5900 -3900
rect 5700 -10150 5750 -3950
rect 5850 -10150 5900 -3950
rect 5700 -10200 5900 -10150
rect -200 -10300 -100 -10200
rect -200 -10350 100 -10300
rect -200 -10400 0 -10350
rect 50 -10400 100 -10350
rect -50 -10450 100 -10400
<< viali >>
rect 450 550 550 2600
rect 2450 550 2550 2600
rect 4450 550 4550 2600
rect 750 -9700 850 -7650
rect 2750 -9700 2850 -7650
rect 4750 -9700 4850 -7650
<< metal1 >>
rect -400 2600 6000 2650
rect -400 550 450 2600
rect 550 550 2450 2600
rect 2550 550 4450 2600
rect 4550 550 6000 2600
rect -400 500 6000 550
rect -400 -7650 6000 -7600
rect -400 -9700 750 -7650
rect 850 -9700 2750 -7650
rect 2850 -9700 4750 -7650
rect 4850 -9700 6000 -7650
rect -400 -9750 6000 -9700
<< labels >>
flabel metal1 -400 -8650 -400 -8650 0 FreeSans 800 0 0 0 GND
port 0 nsew
flabel locali -300 -6900 -300 -6900 0 FreeSans 800 0 0 0 IN
port 1 nsew
flabel metal1 -400 1600 -400 1600 0 FreeSans 800 0 0 0 VDD
port 2 nsew
flabel locali 6050 -3550 6050 -3550 0 FreeSans 800 0 0 0 OUT
port 3 nsew
<< end >>
